//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
cgLuSxoUwnK6A+L1fk12O06CPUysf2I0PED+tJvBzpyKbWaVxPVu/HgWmYYBisfu
pn77IoRysl+Hx9356dvgaL3LrfogjwT1gKPa6Zse3PxhhtiR6dUh4KgbY5lZkIDn
oRffO1f/yhwFOUB66LaBNVMTGCCR+kyVTu5pzk72SzAV2yFZZOVvr3xYmeWfktzQ
x0zbzpE3GbOqlRBeNQLjLOlJqvPw2A1Q8051oNUFMJSFKg8IxasvegUxTU28tB8H
LzZjBZB7VRrPS8xtd0C08BchirQXk3jo2Z7ue9GZfdZhTWAElNloJFblAMSRZbnQ
HvhhnNEgYmClFiBj8NallQ==
//pragma protect end_key_block
//pragma protect digest_block
dZSxjIt2LbUvzh+Va5r2+suVF9o=
//pragma protect end_digest_block
//pragma protect data_block
Z3tcItqt9TFi1ky6Wr7qVhfi5nKguVH5zBQpQNtc4DaHqGWczH+ombGHYRtVDqoN
wWJwPER2NNCEAhkb1YUIn6Xt8muwBZQmDX3qVq1lI3yj9EpxRMHJQl+zT5ClelQN
XaEBw/BS2NsutGkfeoH4xEbBPBgnn/m5Xo8/49wwsZYv2x+WxGnHKya7BKcQ1uwA
RK2LxZ3xTUmDXc2r4zndQZdsk8eGh3iDrJpEGzMpVXTflQ2LmVCOI6TnubdvDBuE
2dPdgSn/6Ic4pu12PFifVL6/Cl8+b3J/QsRfV86OYnuVaT9OcUf2AVVNw8DDaYZq
McoJSchclAmE+KdU1gJBAOGcjXusX0OLKCViHiwwALPpXnmILUjan7wzo3AeZiml
ccfNvRaMM6CTQsmK0z3py2B6X63RrTPrbZ6/GHD+4wX4BTvFu/KJqqwvWHINmVp3
0iY1jBqNU4h0qzply20TJ0ru5kF8q0nlAWuY3h1lDhUMFqtTnjnZytPcFeTJm5vx
bRqLrBLpFRvaohPYvJqPQKwVeUs4QphSL507yfbWuZnuVeN4CVgEu/aFftDThd+L
P7zFl06rL2t8yL1VCDkc9PzPCvzsGmm7X0zdZ0RpYSEaNhK73yioSmgmaJLBIRDC
S4MvTDmlTog4KNIp9Cvr6h0fUO18F4l68MUnmOCS+qd6P37zUGjCCyxkp/Q7UN3w
EOhtPVfUmMIopRIpF7EwbFb0fKHoP7kjLzIGtDywZ77daSUSpGfM4A/TmjmiWYbL
tZflmB0fj6Zszl+N+esnT8abkbjVPgKInAqWHVzAz3lxLgFrjlN5nQ35B1+nIXN+
i4E6NBV/T5XGrbKUjBTfQALmPik/Ccgs+vaGRGVA/KVB6PoS/ynymRcQhTQ5UKA3
icd7gMemTc1Xym9zNXhlxEOwgHxT1xyCg+h47zQ8I4X0J4/C9TJutn1SR9xhkZ3T
UWvBZTMxojDcfwg8llId4jvDR7rOrP+3qHmyeBjFsnIvSA3ybgRbF4dSzTJaEjvo
zJbwKiZuG8boeAJ2yZ/AbxI2oSu7yTRGm3Wx3qnetgmJcJAno17vHN9OOAayp/X5
O7UiVCZjnb39q4W93xvlD/gcvym7dUYWlLFEbZYXXOkB3U5fkwDRe5Dr9ArxHIfd
PrMgu6jYeJx7gbF3dlFKDgwHJhczpzK1wfAcOB8OMNhnOhT/hMlaCZXL47d5h4Ti
h/8jagM1Z4thwXzkJLdRcuW6xaHeEA/lA5FlmpYC7Bxe1YVTRolqipZ1Js9Qr9Ef
TGGPlSL8HomqTPRkEKuLLKklTODPcMHnejekFOXDnLSLe81zi0S3NmznOBxWlzAG
sHhKKxR1/NASlXBK3QjbKYOMTDw+7BpJ25RuTTNyc9KfE6d6hg9urfRyiPqhObE+
5dn9cLrXj8zLTtJbR1Tu/AI3kRiQal89OlzrUPHUQDBoarTVSTbgazWPGSgVWBbg
G70oqsovskmdVPOaCObWUWZElTd93lLXc1efZ37KD5sm6d2i8bAJ+mhJrpOIff5X
avYi5bsj8xvF6idrt1WG6zikcGvPU07MIRgYqNVaUOXGE3gBVQJmQtI0ALlbAOD2
kEDL3c4hg1bJD193MNxGttf6TLh2nJr3hzJyIqcODI0Onxt5FapG1QwRk+yFoHar
0IoodC0okjIurDPJ4MSjq2JntSkkSzVIRvtMtVCn6Vu7uTwmPuzGjxemP2nAjLtG
Q5bwVb0P+z8p8Ju3XRAxnncp0TMmEHgVah3KEeH/IlxbQ+jPOosttEz4gh9z8SKD
YMGZtTEDLCjW2ggvAgDkVZqjEvIU4unTN2kqKZuyS/IEFRugX/3Mv+MB1163ypt7
9/fTYeo/vMx89Fv6wm6EtxNasvQMfLlEvxJBka4sMG4i6fmWjkgneQ2wVnwwZcRC
AnUlRWIxWtETI7fpaNtUYVBnQ3snr/blLlITGMycn9Lv2AQx600yRaOWV0R7R8jJ
6o/cNvRfEDHpwH/hWmqZtiKewwXDBLhsAjHqtISoUIviYl+2N46YSHPHorRh0apo
iL0pPeuhKDKgekwWPQxMcLS8/07GiWp8vnquY5jb5iUIhzX1g/jFJdq0gxSowsZG
Ic37jQdWcymI7D/EZ5qQp450+JncHYLwwj683Z3+3lgiLDzO/yiWMEOPckDb1N5S
3paWRNOriiwjNa4Ju96Y7kNFgplBWRlvSN2i0Q7OyTLjCAcdzMRioy6ch+36XdjZ
nCZphe2TlYdZVKf5cwD1Jmz3GQ9+uAL7rRxWJl9uY7uZ1Z34BNEimmFez9GUerse
dqr999IE2aIfMGiSh3GXTWvi8FYAfPgPY9oTfuf81OPeRL8GuBGlCON2ilzC9NZN
QP6rX5gGAK18ZxDNjTX3T0ld7teaCCQjmt25p5WoZi18RetpT3Xv3WYbph6uk+jc
/sLt5cw8tx4W17NLW9aDo/9AkZW5x1oCQ1H9lCDcCqVmnNV6cxkaaWRTvIGrwDlx
ESLXrbuiF2U2kJ/Yf8ESE1pQpqeem918T9M4CczWh8GYQGZiOZDReyeqIEJWtOkJ
f272yg1MRU8RGY+riCw+KbqMz5dU3ztBDGkg2EFA7VAXuyefRpMuoYcZP6BL2273
5QxeN5/Sr21T5I5fcatHyfAmjkOPPnCrzwRMOhg6zFBB26Q0KEbt+S0+/0E6gjzV
pTh6TefmCDxpt+1FdJ0v3xKAdYIsZ8F7vHvs/rakPWyxY6SFBqrDd4DXKwcnzz25
GJb9F4ZSFWaacw8FE2MIRuUW9UBJ4p/ZKc+dlWwxN1efd0CSlsClkjrTcmsyjfWb
GzolJEA7Gftp8eT5IriERI26XSzDLSPWPrQf/u3T/Ly47lLSNEIwwDHRpFRjBLSr
Zeqb/83vg0LK4nbxNqnOCtv+V5abgbuqf9u/VsVU5cmtCd+bZ0/DXCQeTBu+OSmX
Y+WzNB2zVzIjP+kHnLl+g32G9+WsXUm77K5zGUXcB91NKZmCesCB9cmIxq93BjAg
NvSJoKZTmjh9wkE9VRQn7d08YYP8dWXiFrA5+XgsgNiH5+ZlOJoJ2i1A0PVll4yX
PDqcBbTVHuK0WnKepALUnO6ff1Gv2Objaq/0ifbFXpCdo6XkzBZ227TFcTjvmJ9d
/BWAFB6SQlzuG0533/UmAmintbMXvDivMi3weYDkZJt+oaU8ALVsQ+435Z7MMYDS
tLVh7U0Oo6iEyCL9KyQMXBpuE3Zu38aCBpJ9GYHNORCYl1CHLY9ww1lnCiRv1UAH
bF0+YbUCv3tYFedbdKfMDueHetq/Iw3yC2Gd/FeU6cQw21I6NDctB0TLPV5xqrU2
VFQWUJ0oUoWQ4HEoVUYhMCXh6P+OmFciMgXZfu4yLuPB3p0/Z563ZLqaJAXPmW/V
EbBn4upJLCQQ22SeY12r1Quh//gTvYrPNW1nXOXX5a2JGn0ho9MjXok46CRhSpEc
UmjY6CvpceKNr6TH/o6q7H8fjHj0At8JaewiztPbPif/8s6sDpd7lVge7Khbh/C4
umMVKcZJ9KTwD1ymVAPpTil8dN7EVIemwqBDf7Y+N/G6VrvwaGwVP2Vi6EZDxFf3
RnynA8MjlWzVeLVYMV02dRZMyLzzg/1el/V2YhlTOsozmNEUlvvE1VBNOWWsb/kB
aPXmIryPWnnNRez6BFYrbVF0aMysamICCQ6GZ0wOTxszHFPasa43aQfkvh09L7dB
wHXOXYIIWXZqdrNYXMm87ukoJyS7mKPobDfN/oVHFwuu13jccs8YkoYrAMSFIPnd
gT2z0YsC02RLTA2XoIDhZ1pe4Jlfbi/+AVvDbrnul7XOYLpN0baph9YslMHzZGTM
KnwNsP6wj5FlV5LfLiMWbkSFqRs4RDDEOhQ5zHoraWSstmTBZAD16G6iwz+Mscx9
Qs9ji/1peOVuiTErsWNE/u5Eubbl2xmKeI7QqVmN1NeWdTyn91Q7of5Hy8knPlIU
TmrClqpqv/mNFoVfw+Y/ZP6ECikvsura3h36gw1eWzeHmuVav5GP9LK8bw3zG4ng
fn7WruuO5b1gvkqQRJc/wh9m8XJPlULmvViDrxwFATQE3ZMjdY8TCcHm7HADYXYc
7ubDTVeS857L8H79i4AAMtDYVSNQ6pBa1veKpb2WBQJlERjkReQXJWI4VI6RvtnE
zxkTwby6ifsnSerYf9hjwajqaE23tzovmaAGpWtjlk49hvpSW/Iv6MndEnzHT9tu
FhPlbVsSC2KKtJa+D6NjuHjOlBrE1Z+SeukQDfPI8Q6XxTZ+sQkf7VDfxVchjfjS
+RRkszbdr5KCYN0ZbePSwLKqUs2YCxBtyuBCuMrL1T8N9WSpfs2jRnVH5H+e6v4c
iuOKHcmXQzlxzCAG7hwjTtdlpb+8AZZnDPLDaNtvO3nIp9SvuVIJm+2ZpbAF22Ou
WpeGMKWB6Ie0kxRQze3yFrqk4tFZU1l60IQu9I6ix8oiZwjXRb2XCGKmdHcU8sB0
CZyBRcvFS8tOiXmKiPcxkKEWteOYgx/Ckv4fi+UD/p+uNg8rR1dmn0b+2VDLT9Bo
lpp0C2LfEcVqPg6bVKK8cqRvqnOMAOeWJ4oSwTWb20ApIV9sexAC7e9aRjLOwUtN
kvzHGUYQcpZJe3DHRiTnScC9gP1G7IcEqkK4EOhnvYhgWDVMCeY3GPfWvCgwkth/
nmgpArmjtdjOnqBK3lQvzkjKuFStu8ikTlp5W/onYFl3m58G2Haf2vFCNSMe8+rh
KY0wQ2EdRDPH9OkWx0nkLtGBWZAqMuJva/TtX0TZrJX8XUeTlwI0+mlnRCIo9axH
0hZ5bhMLg3ywX7PijuEHWROUbw5acMmAj7RsZxJd5sJTBRtyPP1BqN4twz//JB2M
WkHwZmoAn9tNpL2yE0C3Iupf8tptke3TH2B2b3rJmIUcPQ9SbpJeANlHlTxeTiUY
ALqaZQQPhfDkhSoZCNsVzPHJ+WUbF9Od+X15zMeNNINP8l5iiXWB3gdcvuK7uS+8
ZpwKczsGRvmnFNd7OKRFUZTXOWniJo2fQRUhx5NZOtRBNu56X0lV4jNbeycJBNO8
e0ckTXbrskHFIwDqRkfzg0mgI+b8rnnVQvw+cKi3xRyTQDGp4ZCroQ2AKJAP4CyJ
cyb3rTa80TsFQqn/LBR7lBWFQRZXCl3DDCLVeFOuvSbIAYBRaua2W2mYxFXUNpgc
UmQL5G3ZVfOld9cCGOPE/xDlPUXIu6Mrmli9RPv2l//FvRAGs12mWZzZDUu7VOnH
J195XCqyZeQWTn+Eyj3Zf+gSmEeX7dawdck7Ef27EitafuGvU+7QRaCnwiro7pCf
lCS/kiDAEg3uB2Nf6PXUEXbJD7IKbmicg1Th5yEwooTY6OrlKO6tuPW6s9xrELPp
0s6dybUUoYjA5ZfRyRWgqxClPzGN+aSCVMD9rPHBPoFTeUMPb8Lnnana/Np1IUIA
8mG0H/Xnzm4W5Srgtlagyhgg37cwQ5AlNZOvs1TJLcmh/fmncOmhoFIOwaLIz/ec
xpIbXBMun2LpeDxV3VcwFU8QHSKMG1Fn8pFDByA9aWCgq7Wtci5RFA8+Z7W5i5f/
GAwSAfQCJRAOX1vkm5fG2vsrapvmMRnmYnyl6OQ/1qkRpwCGPZdcpYtv+MoaHNnQ
3NFXQ16s1bOqJRtarCI2slRANrmEcWfHM/wgB7krhBn/47UgYXF3Wpk+YTTGxeU6
GCHSy9+6cLMP0tLGUz5FWweuWpAz4r1FngrMk+k8GR/FWGzYpMe6Y00dppSa37Eg
bG35vqn2IYVeilhQ6Zs4PWn/6SHoHWM8aaX896uC02WzNGCywOQ/CeetdYF9TxeK
g5qLypknoibSR+P5cyxWNe7BrOmle509AQBm4gsK/jSaCiSuBX2UbWWbER/j13GP
ts+if5T9IpO5cYOIb+Mzo61+YqtkA+nf528RsMWbxsm+OMh1fWQn+RIAO+avn3Po
tMlK/E5fKtW6Be1NJoioDqaT/cx/YZR2Em8SqwMKGEdWb611Rkgk2EMEPkcbQUTu
AWUe2+zADJgH1crE+OynCRcDKTJ+nwp+0ARMhP//X39rZmMQQ12mZvIRXh97d30n
Q7nVhu/asRvx3CFI1eQ7Mh99EIWrFBwRooJnhhslI+a0B2xal42VC0diMe9skA3Q
3Tp57PkFQv066TJEAHFw/aHyHdPlI9UH7Zr3R0E2C5Ex9VHqOS3E0A3bx+kFdR+w
h5aDNcDRANOeLVosJjEuaPqrwI9ivWDfdDq6LS5EqaG1OVjX5PTl1bIcm9xuEgOl
+nucXGK698mZEGNi1E7JFtmMCToflBTrnGFD4KX2vOVfGGhw0o8e8HLWHEZxzRze
jvZiiDahZ/9tlRA0aJC0BKuoQNd8RTGNEnUbQNuRigM2nkNFbTTQ0xoXQ9Z7/wV2
HkO3JrhRbtlYoD3y/+6VIIaSxzm3AuMe1TKWGvA3yOCAEtiiXpznBQgW/tzXmHKU
t5fyTP8bZOeVgcpVrlrlkgkSDbQUL8lxbQZ/ULrKee0YlX+0dNsLJJcd7ZnfAog3
g5/Z5svcuVfkjrcUiFv8lNO2M/oWder9rSLfXSonrOVOXR+LSwH7EG5PP1e2grg3
+MfD7SQ+ZFFpbIxTEZ7LdYEqw8WxqNh0cJXPIiMSoDusFUG9JsApIQws1Ogl0hNk
HaoiS7Y6V3RLhpG1R04uc8V57lcjFtnUv0PdB3f0N02Jvy95fM3cfjKNduDIq4HI
HYKY1cNLdREXT6fTDhOPaPKt5q9VDiODmP7YPuzHtCLk4g7O2phDEHc4EZINK/V8
WBDC8BO12V2+iB7P8mP+ZdYmDsaG8VN3oIKzWNZtIK8cZHfOAodi+GwlTnNoHpE9
Upt7WRS38d4vAMtCrzJQrDzmTQ4jnAOiQseMX9mXfiJNcCmt0ohSDB9BaD59FuWY
F3fVVQeHPPLoHM5oBwU7DkhuiLpii7H3OKYJI+1jRPsfcgLzcrSIzAVeTgFROz7X
LoXF7rypHP9wCHtcArUfaCyXu31jBiEq3t9gZiSaBJLR0W3yxBEo12t5jW2E0vdE
BtR/POF7mP/6vEazhuvY2QQebf6s64pZC9iWE9lH4BsSznddA7vIurh2MzcSjAzc
OiGhXW8xbZniyoHEQEiw01LI6IvEOLBTFzIRrIXfRvFasGlSX+pXw7LHmblzx0CK
wdKJqS93wRh1WFDFtqmAGYzCOBIGauS6jKejGPPpaBtgvOdP5r8b3v8AT8uaVmmX
YuWQH3n7FSFQm1Z2xdiYEel76g9wDOILUfD8b4KMx2tnbjElY+S8sbuWVFA3JXpx
l4aRWe4VGLqx5xg2Z9md6aEWYGfLW+2aq7nSsf0OkDwpOcU5wFYOGOCXUpq3vRCT
EKuLq6BvVw9xArr+9UeNqLBLPlL94GRmySEcTENsz9iQuAl3U9IqyQauglDuamtu
jSQvhFcoh8flqg7pY5bnZz4s6ja2amA6AguEYFpIoakBkJzMNPLTfMh8PIkJZ+3Y
A5xophN1Ai8k4iMNzr8z+bBXZjKVsJJH3WBf2Y9iFDqZQCEhBFqlgn7dBvhNpj66
mx4XOfs/iRVDwm4BcSmFnFHx0PCIObmPRbWOJ6EoYMeReCk6efBdZ7e44qvddReQ
XxxD9GbsIe6MvNxIV/O8bknUuTjclqjaTE8WRLIAXrz4JqKB33dwS9SIkqHfd9VZ
ioJqTRyjUHQZpvY45VkjFZFZu2FBctbCAoewPls4mD+7ts9Za2a5y9eyDv1iAHn+
MzyACojwzcTJgrPQA+ydOxCElZ2Cms7fojeqB4jFYJxoJiQV/nEZ6+jEYZlfcT4B
Ymy7DMmJpBeyhfur5AiloO1VfWLETBP8CHblut4rAFQ3vgV52DOM6m5muZFZQppm
gRrumOVW6oObB/WwkQP3cvn8cHpQh/aE2iJCWCLmiODkKI/rwGGSrI4JyB30GTlk
e2sI9mBWWunoQMjhLC3Hpz1U54z3Sy7aa+qboM5gmjG3l+UHaXGh1cchSn+FSZCq
hI+O/kVN3Q8vspv2A5nHIbtYmmvZrizhAifG+vqSWTJvfgHieWD6fVEUGj+nCtc/
hecF88PqDuRnKcS+VGzOVgptnuv33e/94mZQ/XBSqZDjmBKu/7xuw9vJMs8Um1vb
cQOTrqq2Y6YwE13LqXO4TZclGWcoApUGfO8Ye0GPtwXOQb3JiXCCwVYGCPJ7dvoR
4b/k1Fm065ZBvh1zOZfCIM/l15MMeVb0zJ3sVtSWhRHPfbDd5C1M9k5UbJ9emeaC
I1+3VcicYpo6r4XQl4Sg/yPeaVXHIrfEWii5Hvw3yFH+g23PZ/ZHmL2sXh8RCBa0
ca+C0xqeGQGQM8J80bIWkNmcFFJZ4suLntvB+3wvQCnLOrRmNK8u4XA+X0Y2V4b3
kzbehbiodsZ6R9vFB6eThVvxXDhBIfLwnQv5O6EE6l4KhVxycOsD/2I+juR3Jb9l
CVwKUhxUBKXhO+qXksaNODv1I59ITVDJEZv8JBdp7VbLyUlBmtL/vCVeWbIkI0G7
BHzJEnytWvqadqd0l0JL/VliXWEE3DC+B0sv6nV2TuANnqodj/AwmMBe4GNq1jES
jZyhmp+m5Fy2wl4txujaD/xqN8qUMGP732INUqgME6LX21sl2XvT+5MLS4cjVF3F
hJcjGIfst+ewtzB+obnSJwf0N4uzTLUukNBmuKUlJGmqermE7zhSZHBIgjfsQcKb
Gfrr4pC7LCYogYoYO/o+z6F2J06dgp++2Mtwn7QfD7boRG7L5AeuUNRQb1Zih6JQ
Y6oeAKMNlMYTfL3D0tI7DPx4LzI2cmxRtDTGSoH3VzhlHIaia4W3qFhdrT7LYVDj
qptkAV80N4yyxEdnrb2IodM7juTSIpKkiqpsXPJoheyYsaukxVofn6AIU36BhF1w
rQZlyEwi5nnAp6d1h9PhOP8bTWYPMxf/eIZ9rttKxvc62t7vxSJ540KzUm9iVByu
bBaKIiwXd1hJmfL3t8Hn9okzkGM2adfB172iHxhWoAMvAWARoW0riLC/eT9XFi5u
BlDS3U8y7Tpe0Phcef50tK0MfO257CeyDVk0oSWr01nMSh+18vZl4s+FyY6aHF3e
mLrWLO2Euax2GI4UZIdmV6+uoUEWDNkww5yuVDFMsNkvjUcU1FASE2vdbaMk97Np
Z8KaAiLHFf4JvxmpaNma2DGsKD0lBi7X2KjI+0Nemw47hNirzFYj/zMXODgFZMCd
2iv+zDGxireEF9liCJjrkVXqKkEo5H0KKKk+d7nwqwGzfBEi7XnmsQ+rLNzZYMRQ
DdJsAa1eHOgfOtcUwLrmv0OSC1A7leo9ax/w+VFngeFz1VyMUHDiH4UQP3vSEocJ
rjuS7pFtMgHm0Oy74KmQcjHhvJwdfG5Eu3X4hXUoaWW7CKRYHZr1MEMi14HO68ho
c4lrR/NeVFjfvRBwvAkqFjErB8yBadku51wW4oL/7tbnpELAYBWoKfgNcgI7yNho
OJ9SeKJL8mM4hW+9zOlUxeGiyAA3ljcdbnv1uzk7QTpzeY+semIRagl7Tb0GpCDZ
XEpqPBdZ7dM+MC8MXSdy5gbEHHpLOYEK9dLJJq8LPZuHo5nN6k0QLSWde8rwn3KY
8CJ4625kbsfCsnv1sIX+sjYqXFRFP5e8Izm+ccDfgSAB+7AEmpSK2QiB1OTVgf2C
Zwyx3YJQBv00lI70bvEuR2O0Uio42uQeTIoTiKa/gEHvIVZjuf2ewylkBe7US4Ix
egdnF4Grz6GZDufMJ/D6AzB+6FqivQD5TXpqsm62WmsfYlib7utcrQOJbFoPZJZ/
6etVOpDwnlYdBhIjlMjhZv+ucrIIKrKfp6jR77LlLLhY/ZviysTBBgnnQV1IJITQ
NXI0yWBldGhJhzf6Vd82I0MaWVKdfOWHtZN4VQ0p95DRqyiixJTrNmA1v4HTJIZV
H+GrtFQ+t2irHcWEFw5Lg7C4o3GYNi8nXcuhFnzGqUPtSMIrQWNu0NVsFZGD3YTY
Cr6SIjQTnkC9mZS4VyEP2GsVgpHTBTPou16+NdEp5HYNo2DPR57+pU7DXt2nSMrM
1Bezo9AjaPawwBsFhpsqqXm77hsGIq/0TNIaTqE2T6VtQwqdda9W3QpefcIRVmSr
m6zvuIuvIvo2+1pOQ4RtlFKzaNji1cKlC7VpCFwQIqiql24wvAoU5mG/JDXv85Bm
GGV0RV7ud6OrSWmtXUhm0z8TKmfV27MzOZlbIQb3IPHcQH/cvsKg4W+DBrBbSYs4
DbVjZRlabhXhvVxaXpiQTgwOj0kdFvIUpyTL95rhw2E+0ycyxMgIHGGVMC7dZrvB
M3BDWi8cp9Wizh71ylj+cbEA9pdEGElo0Q27Q3aYMlwYMYlaus3azhenw3/vtwub
7CmJyGm7yMaaSwx81znRTsHxXtJyyvzE4J4PXuZ+flVRHSstSabvXKuZGQgiTwc5
PIUzmow8xllXDgKLqtb+SKrtVWFHJHhGp3I1H1/ZcbC86sdyaKxWRI8KU9ExqLcb
+p1ZWjWv5UaLaWG9cv/KOe6yCxxXco16m699lBgi8u3KE+ZlRAVOVqJRdWCgXB7l
SSHWjkX6T6UOfuBAilQBuJnAX6Amk73kJVIbgm6dMZ1g2Mwl4llODSeh1344jbLA
pVf0F5PfzzBvgnLzlETVcveNVoS634jBBfOjFJYzEFN3KM5rGiQ/x81RgZIjtQ2J
77az+FtKdkV60L2JV7rzTlrnY5XuJDWTP1ROFSkUBhY8DoeWh1/FklOdjTeAct7h
8HwaNwto492E/FsP/hMeBYpO8ppgabgXwo/pNgoSBmuQ6hk5sM7riIRoadU56Ngz
PETfjqPkndctlbV6pkrPIPHg75FRiS4wXGioGEwZ7jfrSO2rDcQlbhOmjTCsOJ3/
YbpIcGb0UvO1xPynhjO4YVdTMENkIGZxCtEx5FoHFm60xBPWVG9hDhanPytvtKva
Rzcl8gGX0qO+EQRnowlTWcZaIThhFpRxcxL5HwsyT6nOj93Bzpyk7uBtg+mihe/I
elMgjSl5+edyjWj+eZsOTTWaTcp6/0IdZklaM5cDxLGka2c1FEF2r705CGFU6iNu
Uyf5UwQxpxYvNlVCN9gYuselqvQyX5d1V/RoR3sUQJu+30wL07BP+xSV0Zt/ASuF
dj324NAHtq4RDmQfooLQvUPZyzd8xtO/MxUQ3CiznHltwEYTi6o/gJhBXldslnwS
qcsl80eR6AzgLv4ukVHEXHgQzJbv4RxeUbH7nLl6X1NXWSXmRR+r2ciKYjsjPzfb
G8RC/LJNHl+Q9ej+7k6Nsg+GirB2zIgwa1JmuoIJCMt9LrrsC8h96lSHwWLqkfDl
FH+/sT4sSJ4mi9IYigPMHkoHfseaSamX5V6XZ0ANzjf6nRb3kirwI0HxTFUtTVdH
yF7vAi3276/wbDyzgo9NYWqG+QIqVJlaeenSWOYLrwR4razp5RWPs6uqYNxJz5g1
H38BI811KeTZXGR5oGn5tDIBXePLAgZ1gaVDkMHbj9AX0I7U8sHpDe2COTEoI3w4
9EG886ydiqdhqLEF+hulhKRT39NH/2wA3dcW3lSnJpDsIXmNQJTyAP3uVCxqT/45
pHqywmOwb+iVXD4ypDn2cUgoG1nbOH30OWIPQqiClshgMDl/7CAj1qaUJ5gObow2
pWTee54Vdhz4NiMkvjh/G9j4zfAr/c58z5sP3hKSsJitd1rSdZgBLXudJQlDpnHJ
vgM0oloXxd2BriOpRNRkyNiBaVB+EuRf3UC1suRwuHHYEsJE34HvT7CPn3KqmYbQ
1Rn0gu189j2wyf2BFM3vqE6QJrwf8qoklztzcOvUN5FLZE/QviiIXnqA11fHWjBU
kqUGCn+tTLNiPJ7CGHRnuZ5UsNmux7bAGPAEKyojTXyUywV+LDsFRnw2a4yjakcL
3b5X2ilT5RTIL2BOo1s8O9q+0KyMvLBQSGyvkmneU4CVmPXXeoWm8a6KIpEXdGko
VHcVKdWjk/cpwLzxRyoWeqfSJq7sDv5qzjFPukDofjzyJA8IkwHPMwbIvMN4PYQi
sz+/TMI0GSeePbx9kKw/CjuR+UJ88z9oPRpNLk3XzUH/JocjQm5qi1VSNFWALwXq
6k+1t4J7lcqV7QxXygSXT9tFEDXb73/+s6h9BAuujuE7ohNhiFLn9Y7qqxH2iZnJ
cvebfUDDwtwXXKu/zdgB7vuXmhJ24LTe6Y2NZc6H34WxJyK+lKV9FQhx3vczkXUD
ME4FjSsEoY6OaxydAeYlmguR5UqlLsp3c3v3QQ8SctajCTCmmFWhcYgsoSOXh/Lq
sxp6vr1FBXWWQT/HEAanPd9MEq+pSF8siD0ME7fKtW2kkSG4el57XTk+02hBhkAs
u7cx9W/7XY/Ck0bb5CCM1qsX4SsR5aXK4tTZVrNtvInKYsiHQTiZDrcaY8SS24Fi
wIFxkYa/sJaUgYF8AHnGE//Y12zi025Aiw9w9N0dlXzdExvSTHbtJOaz+CtfKIy1
iGbJls5kEdM/ZOqeW/RK0D9RAfkasdin8sVrzoUuc7IRZrXeWDQMAjTXkmP8qiuK
rkVx+cHcNXdOcO1LQRQ/liMNz1Eii+P5JKIZNOZEEf/nbs4DJqaDxhTIjC12UFra
IyJSKR0hAX8K9Y/Jrgt7abIKzXnw9w9wRTTmk8fO9fImOHcB6HJgpwOEoAAu6z/Z
gjH06CXsEJvuP8sobRAug/58Cz3LrJ50rAuDlPJPav/0nN1GPztL5Q3XEI/UtgVD
TEnNcU5dwYB6pHjYsT30NgRohgvazIfxGpgNqnlRoKq8uQuAfx17HWSiBr23W/uj
0GVzZdwVJRX4T2aOIdFZanJffssud9v3Dbl7DrW0jomcXflDAQppF5N+sHji+Fte
5/A/ASY23A8KMQHmGjdmXLaOtkcbSZCZS8Hi/ZbAKMO+Q8aof2kAcWSTkHObN9wH
9h0pCCSkhG7JGzqmnzejWgb7aWjgS3p4DNa1s4NEaPtekwge3bNqESFHxFsyg71c
JAKQMqLCAYO+saQw4iy9AEpuMDTHBDAjLamSk1ZlD7hFfi47oPSOPrNL40km/KlT
Gu3GeJUB7d5DYvy4z5r2C6W1yJG2iwG68h3zytQ2Ncxugbwg/yj/w0z6vsztQuiO
GRV4ktToVmwXfnT6kGpqAz7k0A43CAGoAEDinNvrupRzVrdG96r+U9X+V8G47sa3
48smlYIWewF4JKWD4azkXPJTShJcfyxCzrDxj0vhs+zhJEfn7icXAJYEl7SxxWIN
lgIG4ufRtm0ErxE3zUGj84kA0BTgbyANXciuqD5ZG+C70T0icl/w9L+oWZWtqwtA
Ai5GVMoG+nT5SlkYtta4ZsBKGKTkvMPYgyo7YFhYC9pJn9l8AM1bVu8+YmojwEI7
aplZpAqUl0wdMsb4SeX/EUP4TLGaxt+bejbd54EFd3QlwRK46jiLtldmLJpbh1Ob
ny3UNgSzC2bP6287GO5yQkNymUTeWnH9SXfZrNQP4+/bt54OqpdS89g3FwNyGo+N
aVB8GN7862LngUh/6ci+dPGVlk92v4Tp5ImDSMC+SG4fNVIUviVkD5NoPpROEyJy
fBe7FbSYoOzwtMBZNgX1AfGMUiPIOsJHB5YLKKXjaR/nx5M1+8F50nQ7d6Rrgbbv
uFv3e8G8RlVIqRedUn/eUSQkYUH6d/EVlp5c3OXjrTJnXpmmQQj5KCVtBrV4BcwW
y1nu9BG5EYEJs401YejPmBolDoHJAU1DQiv1+/vp3xalMMVHqj9xfioL6wCOp7Pm
aAeGKRIsup6gxpOn6+peksXIRRWS6M58CaJ0zwKY3KkNNs1HSmemkKGBCrSFtXLt
JrS1giqEu0HM7hbwdyRHSy9dLRej2vXlH8FYdyChpaQ2tkee6shGz610C7OQP2Eh
VaYi3cIg2rIwNPOpJhpaeG7UiyJZ08mVv49iBr28jgy5eVMzsuRZ1vlvNrZBWICs
gfsMiB4tUVbJ5F140Leypv0AFgx3G84IVH8PxsurVuRRgQkaiL2O+wVskUNKMM02
LLLQQtY7hAhjtlKjIavZjmpALWOMwuDQ7dL98mPBi2/k3zQx4ZA0blUPpSB9si0u
WZP1OlQCmkhchirhkZQ9opsUHg/qPLlURSJDixOd64zcZpOSlFIU+ATtzwQ9X0WQ
t+pfKafPMeSH6QhQg84/vNgpuZw8CSFXfmFr1wXnS4o7MsWR9vgrD3hsbOFdHQZf
TLxLCkcTyCiqlqEluZZvpfNiRxfrBsAlOybTStOw514KT3peTqOuD/qUj43SXkBS
kKqQi4Or33+U7mXG5h45burHq0aNZmEvcEPwANTVudxENtpTP0Mn9w5FliNcis+M
63jTiCxGAV1D3pUizYp6ML6uw6lCx6G+gJDh9JXLROkRVdeZzOpj1uTUcPWFZNui
Mr8sole+eaw+TjOiUp/AvvLRcMNBPDpOPqN4qN9P68ov48nT5pbzdhAmH+HzDP1v
w1z/cBN0PzfFY5dU9HQkY2hmFn/SsJajSyO03a1jpBElxqSjTxPjU2PeYHR0R7dh
Tjk7PpXwVFAChrteuvVU1gg7Qp3opkkOAxq1Zy/MOZYDKm5ADlGkcfoDeaDfrGT0
sZ9ZT23oA7mYrraARg3DVIOs9kO4SVkXWTD+wkeA9J+8inOTw+bYgMDqTwW3Kj83
OePWiXFr2Lg+phSQb+C4M1doqBp/JrnvB0gOa6j93oZ6Bsknyl8WM0fNOR2bxSuA
LFDGBYzOp/bK4fB6EcyoFE09ue3Je4F7e+bBegH07yA2X2UhhjpCMwZYb2sJDkC9
ENqOXdl+4t5mzJ6h8TrM6C7SFGnSFATk0qFdR4BBDcZFW0FIce3xMrttTt0zYT2E
LTXHT+/rhqMi86WL0b4rpfwl35EEMsDHQYGj8OHBpa+XwTtrYz7Ia3s/vPX+1V/g
mChXQK85bSN/wBseCo05byPb91bWjZbXPmILJLC3Z7LZs/WeXLcbFiJJ+kobWObw
zh3Ax4R8QQuLdYkg0s2l/LPIq+Dl62plbSoUumZmWr/nvhHd14orXGQ4jsYJY2po
ixuThIO6yCFnr+5GUheHmDFxpn3DYmZ8ZI1ArRumvWxGPtfHGQBYr44clQknM56p
A/vG/vXfD3u8gvKPsJ4dbC+eJNw1qrkycwfIb21swCrlBd7PmTx+yzcEXx7Q+m93
vgR4gtD9SMiQHN43UrasYQO++kUcEf74aQqahmc+R3ZwBBlWRdJjSpNGZofh/dU+
d8ZARA7jSn8GGK9dafcuNMtFJDZs+yxwbUF1Hp0pMviaVhdZXHedDvuKBI5O9PPg
KM2Fl7wRqLU2BFiGDRP52IwdrUNB/qAQ/2mYSTSakMgRc1ibdij0xDdC4BwlcXwN
7AxJQW3cGoSzDbVfgP4u88mCdk9AaZgH+mTJFc1SJCZg/+k+Qwh7ORxpbfofIt2M
BcOw0siqF0ESjmv0VDdyRjGZU+zuiPukP8bRudvvE/A8suDM95KiktnKGyLfGPtY
q1vM3Oe6TOf1wOCkK4ZGq7/ZlweWXJ7GX88HiSDQfUmiG/qfenghCnFMPjGnFUzr
RI/rwIGNGoysWtJKJnlRNh7YMKtPCrpqwYeYNrJOoHKou2PPzFoC7tefpkK0kpev
02t6c0E88TcSbv9GDBXlrl1wxd0pz3zExIrHLPi+VBRIrFAx4ufQQIPP1Sb58TIj
e0PJyJewtU1o/bQbOUSyVIqAKtGg8GX4NnnvryizyaFFqUe0m2pRgRQyB8z79hQb
GclrXHlAaNYp+De5TvsFoAM3QKSCnsIS11do/i9HYD7z8tlGPBDxsJMJabqyen+o
2fn3OdaZt1X7LHbR5TC19nGdncSbTq1+ZSeys+ZsjcAOjmI6tuapUKkWGTwxLNu4
kkWs7Htg1bq32aF24F/SJDofIx50JgVboWAHKSGrHaierZNT6IK+oVII6DzLcwRW
6hJS2yY7qKZQTItJ18CLVYRViqjr0dyCs9qfuPJUigNZpaSpvSc00/y1y3tpBlJV
59lej3n6WxtzSbLjmtt9gKQT13T+WJkNWKuMrlIofPoSr3XeOQjWOpCBvvxX/Q7o
NHSafkpLoHodMjCkMJFwgNzJsD7ARLBj41PLfDAJHUxteL1XLW9g/sFofXr9vTKY
pvuAoMRCKI4DUf9NwTq19CAMwf7qyliwRMsPg/1yhhfum5PjvC1SUC8NDD+rrDf4
24vaj7v+V4dtUcdSPkCljoP8kcsTXblh6mHNOTIiOdK7OF43Yu+QcXYz0akmxrJk
60W1JtV7iclRu1idL9JNYL0Ff1NVB1t3idSHdn/iJvkIpmhEh6+5MtHaR2rQCnIn
lXCyqVje+M+enjeOYRdickMd+pq5siy0i3qe8UR9AHcOKsWDcxfEbyWFFc6hCrDt
txDXdAg8lm5gcHfbNS2rdtfetB97w4MzOSOTdk9v7cJlLzLCvJwDxyxKmR6ZH4lG
TRg4SUNTHVlVUmptBYrORcg+gH3o1MoFk8uL6BXz5jQ5s2J4QgtDGsyGMBTMKAKP
Y7Zw9c0gOXVaVOsuwo8Spl4I7L7CEioo1DLLc37jWCB8+vndiMG5MKhpGMmyCeYJ
VpZEPofYijvAbR+V138vszaWgPwKnw57TJAdEAhVz+r5Ww0UWj4sd+1hISyaW86I
kmZGVNDF4nFaCINTmdkpf35yoNQvnAtcTgc0UpI44o3FiTB1By6RFLvpZ7dXcQnv
w03h7bBQS1lL0YuUbbVVPZhX23YpPOXX7dk27Zydr6Y4ZsZsE7tbW9fxxQmJJnCq
ngd6qKKoAjjDU8QkAxPrmsmKanMF0p7iBTijHld3KPGz/ph4dnsZxAH2a9neL9HW
GD8FFLtiAnZV9jFRd+Jf8KzpdhtwjC8s6z4Abmx55ejZS8SDGLoL6SGUl83rP2d0
JuUDwEYV6jq+jJaTWwWK0UFiDn1OHjbDwO3Ry9Sm/fHfAygSFBuJcaR27nXo0vJx
BPEhhptHoWSspIj08LfVrc2r+9vH/6dncDCKgClpRwIxWmbG85mpqN+lqGZQo827
mCxIZPV+nYL9IUdOJkBTp9VS9JM06xt7nZ15U5xYwxsnZyJV2KC7cF8tgohRKUY8
/kenZ5cXQ58ACSlvlMb5DwUuD7d8Frb/ahfLGw/Qj37nDBvCXMV9q7/yVCgGWrXs
AJyJ/FRDmz2B2rLnAWHLMoKwPHkbOWS01SjNQkHshA0m4dzIRUoPDI2WLzMPMYRa
xO2gwsQQPV8EOuG+HXXNzpdNaPXF+TBMnNuR+Fz/EhQAaGXM9YazjcWUywy7oWz2
SrM6/+dcEdDEM0A+Baad+eFPpSPHGJORKcc02Rg6Ds8mFuXaWqTEgLKgweOaIpgG
loQFjula4KBVSjmDVmuC+D2LeAR9Y9NxF0g0jh3SnheUStPE/n1+z8NBL+wZpUsK
BgEmQ1i/6Ov4y5sJfuCD8pCZ83W0xFebe9JgjzgVv7U8OB0MMTHzs041hG1NYbPP
5DtPyk9ZCZwsYmQcF2txv5preGW/1s431Kd2NbCW8e61xV8m+A9eZ40k0IXfB6Un
2aNriPaNnL1JQwQrxTvWSfT6xr2h+qGTlqFuC6NAgxBrxBGlplw7Nmec3Akfp5kk
/eShJpniW3/uqQbZlVkz6pDuU23D9L2RWc7OhPQMjBXhI2lQzinic7ytF1EmG2Kl
FsB/NxrDSV153iOqAzHwSZxkcYHMTAdJloHlfwwJO2QLUxJItYLunLv6aPva074j
Aw1ZQkGAqAixAjbtIngOcCZH7BCdY+aEopK9KnslQtxJq/lxulb4rWIX+JFhvLh3
RLO37MiZ0rNi2TQwPYbrxdAY5TK8RI8hhfPbdSM8VLyRoEEXJIkxK1z310akU73p
9vasLtNbbDqNDVuuTYu4hI1bdTgmTpJ5xwmdDC7jUerALpQxE+lmgljAcG7FbuB1
il9hKZI9fXZdine0lud5vF/S7Hrr8OJo/ULykzAth/6ZwxT9ewlclQo0E7cnO1wW
4yYwnMhoWFKKAcOT8RteXKTe1weY/PNS8mYKmVWHS0BFlmKz3WZctQ3Kv8iPwg7k
5kqr/ALhrASsKgUdhh0X+L9EAIEeTj7hQbGx7+dkXDOQD6k9ZS9asqwl7xI2iKXg
IHtN6EEhhVnwBraJpDma00A5sfqdy8nOcSNg+FU80EZMtgBTgMD6/VmTJ2XxIi3O
HqLjmKstgizkoZGV2tM84X5TFAZYm4HufX8wudqRBnyW21PO7iQYf5SGGAvBqUS+
LL0lDU4jIESZK2Ao0qULH/ZMNSR/Qi7/iELHYg+k2WA7pnuFZn6c8zMxKRiG/QjP
TPQxeaQ2l1QBf2orKFC/gZzeZYe1UE/pPl1S4Icm0qvDExPGrJVcO4U2CGBhHdQY
rzW4NMtFsZbzVkbDZgGE2+3UvItAcYDOuT47WTde1g+JpkElciOu8zvLhgot7pm2
fEz5u8Eo5TrcDSBZ1sz8Ru4L3ZJkdIHT/HmdUB5Pt2/hPr8iNQsCfw5HO1oekuxy
QSg49AugsF2VBJxfn6IhQAE+5Cv6h2n6uzTTDduOFdReMo+NA28lEvoD5x2o9E4I
PbXpPRKhNYftmD24baOOGw6xELw3ACoq3xxcFrsXq4f+mQIYyLtfzx8W/d4k4EAC
ObIpI5e21foYvmXhpnOvy4eWutCqZt6sNRwAR6/QssHRkeXRP9IIDEZBqZ1IvzIJ
ZpsBHCqT+tA9vVAsiL7yNvSngS2N51cBvEexrFD5CRjKKiS4smlP1Knv6+hvYGvn
8sCtF8iX6A/JtxNmtrMsxe0ToxA/PDhcIaBYB+RKz0GmXqQEiD6EKaOGuVfiGq29
1X3ap5qK7VtFk4e3MvtLolY+qXMAVlS+lSL5tkPkY1iCtCaMwlbrdkHUZzjeN/rv
ul5/jp1XKPMejffqMwkGdDSdwTmh/1dZA2WAWxxfvvClbzTsdojMcNPZqG2yPywP
dCeJkOLfMS/OcM2/YUQF5u11szFDjUzaO9iF8n85qJBFVgZyP0izg0vitkRIy6Db
2qbWYD1/O82MDYA/WdDvW6Y7up21p3JzmIXQYqpvPpsE5Gt49U35J0GRgBqe8rm/
dbyzVBxjn+LFL6KCeECLafTT/MDU2QSGSCMc29NmH6VSxgN/MfRFbsSvO2yIWmr+
dhz+J6opwKXKtDYZdiedmIC+xhgeIDy729VRb8nEtJnTfBSg7ief6SbYc8LDsa3p
5iNsm8yJgyvFPkWi8fS8JlExRDPpF97qsrN6qfCm1F7JsKhl5jXzl1eb5+Ck3D6M
cPr1nECz6ZTGy+UpTjRxGDSmkk9cnlvX/r9mBUC5BuPdy2HMTp1732SYLeDT2Roj
cSwdDEftyUOGSd3rTlhXqpV07HXvPLFUjq/LLVMKhyZp91Fr1gdMPN29GMHjXpwm
EIOlFkMQx/AIv6zZYVsy+XNDM7c7H1XsZz0SSndipP6TedYZJJ29H27P3K9ah3uo
cbDWBz6ga2y4rGHZeoMS4f0PokWwbdoAvy3DvQv6THX4Z+OztHrJ7l5TvqBk6trK
3zqoFsPjw4yt/S6hRC7Os+Ty4qUXPTCbkVz2D9/3vGVDd4JkWbOJ9ZC9m/zqgwHa
ZeCqreHgz5bbA8qWmOYX7q6yyzTTRQ9gcbPzjjQheMSNsXpq6VZvgxgfDt8DuuFh
QflyIPU7t/Dbe7/MDAxIEjtff4ev4v5ge3akgDTd6L8KogIe6QnghyNKxSBRPNlr
m/SGiYuXt1TPzM6Ng/wnJ8pW6qFMVP1bdqyOGL63tv1cE7dq+YmbdkRvGO4YY/hk
gyk3B03Qi8UJtFJGbbJatCEc0jdEaUHKUjAL4BW/8mJeJdaJqau/tZxsi4feaBkW
T0SKSmtjGyKt+/aE+qTWRNeXAoFRia1oc9qEpK7E+8DjpzS6bgNb9mDiyrpHUXgg
MsglzH5yZRDuyAa0ptfcqnVJjraD3nzSGlNltAGGXRPt2FwrVJFkjsL7yyHp+Rc0
evIDSIvM2FacYzolyUQcmXrgFjbKIaI44SZe+9T8QaELwTmAvFdIGWWzkZm+2DEh
XkzP1pl3HVNUjBXIoRAKBayL3r486T0usd1+eZXVIYXQs9TM0T9PYBGKjgoJmhfq
yI4OYNkDBztx0UhsuT/mK+z8P4VH1SLkH/7GzcKfOhckl2AfaV06fueNlnxCUB+O
DTf4b68q+7RUDxnHEyqcFmeQNcM8lb5czDGu0Z8R3yH+7OVBpuDklImvAQoQ1iqw
M0nhABpJGXvle5e+rOxg5qA7GC4b3riACwXeXJELjnN3SDmTiTxaSwCK8mkgdSgX
v6ksK9EeI3QXlOexkMfv4IM0GdZUboGBWfkUQkyf1eguCk28tWOcO4VBpT9SNK30
G0HSjUheihZ7tcOgBnPmz9Y32ajuygPFc7qykFUlOyNK4X9hM2G/Z9kKFACCyQyL
xxeFA8yQijKk4u5WC7HbyerbFnGRs4LWSA6oXkBltxl5QvuaPCiNSyrJgp/oISA4
3Sx+vTG+rKZnWYHqUElWI+QqojQ4Nm0OABF/BTqBKItlYVj37BaIAjqFaAA2vtdC
qRzJLkwFmL6LgYX7gQxf8QKisqGpiCgS3XmVtaofJjWO2dJUckSC6lSGN8XJU3eU
3TFAm3oElsWi2/41cjidg0Bi+bKpoBG2PHqSwhBb30ZS4mdJ0Ng9bznleSvXVOnw
THhEPvwRoXLEKnaXRd33rKwLnEQiS8mU8eeG9AJPqLoo2FCdSHUK2P7qrmNbxYO8
yzb4vEOTkOa/XTomwafZ1sreEA9qsoriL9aG+Frt7uwZtQmJ9iwVaqeMQEcyRVFJ
NWnodA8z/jWWhjMxJVCMUhLQv63IMm2Ga6f++YJEwaq8Ep72QRQC4nS6I+K/yN8v
wttDWyYX/ZyawLsvenOZ4DPDjDsap4qF0gttAYgTI9z9sHDHJV0BkUlK10Xdz1SH
wiYC2eo1bVU8Gg1dzFA1DBj1hP9EZJPU2kYlfmQsYXIlGZuuE+VeXkyHo79eABoD
gkOZnH56XlKtHhRX60rtFwofr66AcQyrZjkYjkVggptvciULj/gCFApUW+xuZmWO
EsRhYxvdArPDSkc3N5HAUGAhwdjK/9A9CCYqf/PDdVjk1NYXMLEMCvMPv7vVYC4y
ijBC7v5wzPI2Xz30Z1NMcsqBpXAo85WWtaERZgETYtUxazTEvuANsohFqTF4BtgG
L10TopFn6Ez0armVzOJkdiov2Gn1aRci1UHRLMvnNU7sBoGXlIooGFABuQ1VKrT0
aL8dzTzKpWubFePzp8j/iRVdY+Ag5aPkEKgiWxkDtHTFunhLh2hck3LNTl4hWIU9
NLpQgyWXzhJ7YCr9TKce2k55gW/7jGZPikQFhKmLGvI1QcoT03SVh705RngxSEoS
Yd4S0KHFB7U8gb7Rxhl9c9RGKuc5U2PL4zayIGtDdbFM/MJYCXzyrdMwJ7ri72uK
QuAsVGTbxt44kAtQWChDDA4AsjK32UseKV/hptWvFtII2yGamLbrYbPw8kPOi3QQ
4VOByS71YF43KOaeXEWWHXjYs9j91WtxMTJXXD4PUcbmUVGWYRIaucDr9CcNOdWV
H2Yx+G9+E8zu6ribykpyKn6yxf6e76do9kdy/qYRrSvSHaMTcIJSrgWoZxzYxAD+
nxBQ7IVkwvwI4NfXKJjF8laXlAenbFu+naUbWTI2gyxWUTIKb02iWI+zSqK4xEss
2zLh7mUvuZs8weepEjMFuqRDqxeycndDi9IfG1NU12y9jddrfpVSUYj0lU9y3QD4
osAd7tOZKqi0vjo5PF8/NqZqxANjjhDekfVbseM+M+Go7PNspNsxLFEB+otQJAT3
7Y0OWZGhO39Xlj6MmHwKni3Y0+jm6/yiZ2+70BkdJha/CgrgiXi/P05ff+M+lsz0
BCHGpZblQpDW1VGg+1ojgW9L4HtglQoO3xmYLFnLeB85tDxTD1HsBQ0ICiesAhNc
ZWL2bpZYPLRQep9Xdn389KEXpPOFvpVLNhyxryfBKLs41FGXtMGBwgRDk2LFwuf0
lCzbxmV4egzZ9UnItPGlxBy8dEBl7ccjc96Zl3e1fMq/MM0zTheo0VZpWTRC1xuD
fqKbNyiNmwe5+v8NQCSb6ppMQkwbOS/JOeJttER8FhSROUDe8n+wSaS4C8f/kmM7
8mBwmPfTeYI671GCr3JN+qAfRMG1YIqAJWRRltazreaWSfUYfWNRyOqSELINXsvl
BTpFKZALXfobRS0nZ5Upz+j5DGMpLVis+mcNCP2eu9v/Cc/4Wb1H1sIgb0X8RLuS
1CeY4wKL3HqPJkU0trQHXh/744C2CkQR1mItPjHB54rt7UYCqzeSEXl+gXL16+ux
w2eEzgpIh/OoHEvJpBC4r/LwqLVCPN5LWJIwh9PqTTYn3cDZgKEKIzaCDz+bFSEg
TWlym8ocjKalTw4szXWVE6NhHoUGPXmL9uphFHJ6zemNvmX0xtQDnNzfvFYQwBrB
twwqLmU73urpqRQA+sOpuNJzjJc9d9Zg4YInwVw9quAbVqIMRXFgSdAtnHFBjbvM
zvAn01hBsKePeOmWdOx2DvgnKdPmel4ItH/5ZtajTZXYyavBxZjKKch/HEk5A8+8
7uyeKQiIfYVSsvZxtf3dsGhc2nfDlIWs9m4LPgUBqiIVXvW90tRMnLnoB7jKIcfW
UzhXCupoMcYbZg3tgeUnDgPGaGSxkP0mcCmgogmGLQArytxabrR/RTewtuk87gjb
9FJ9F06DrKaYJwL3+qZkGhS0gL2OX4UE61l5i+pagrSbmZ9ZztpfdB497ohamTAh
YX7w5/VEnFUNCx13zm4eBbzBKbCqsXTXuiZD0JSUGriiWT84da87rqn1RnDyH0eF
hvyDy+V97FpYDQnkEeWfwel0USPu3YaqhqpgkCxLcvAiNR9qCLg1J39/58D1NTHd
8pg/8x6unMuXdFMI7eZHokncuy7dd5vHPNdCPxc1i+VCy+7BKsGnNgM1LSr30Gu5
0hx1wAwZl/lgXtkANNdo84j3fBuDocI0RlT6YTpMKI88nYDX9s30pGewraGyvCuC
U/uYA8esIWbVNibmfYNIJO8rHQdgj+vi8oFCxjCRL1XzJ3AZw+ezO/YNW/AcvXqC
uujMjFF2Cx6ucoE6goAbmUsBbL0FqsAkFH6m67rg+DG/d4VZEFaUboYGaH0FfJ0S
3SKyjraZmC1MB1b+xRFhx1fEa24m3lksm53W+E6ac96PpO3PX6eDkOANSTc/8E50
J+99QK2Rej11uUTpZnsSxChiZylsT2qG5m+VoojQXl4VsECxiAAK4K5yutdUJ52U
JK6rw7ytfBPuWntO/QDB0hNoMYWICHxaSJY2GuUUOoS+eTudwCosnOeCLrYDwRAt
FiTWOpZfIbjBxpjPmktQuCC20WE7a6kGC1bo4MqxULpH6qbYH7TPuMrRQZsSoLP7
gK6IbpX01/fG+zPsr8qESVJWOhX8u2qg6omNA0EZ2tPZ0tP5K7QVI6tBvqz5JArQ
Z38O+G86mvayvv3nY6jfpMMe37e4e5Wm2AjrbKkbc4ICG3z4m9nD+Dc3wGViFasr
jfoAUZ116aJWlB58L49S15RMhbqrdIhBXhcSYY3YFWUOigXX220PJRm+9rv+prBN
PAxj6K2JFqlyWAzIr0knPAPnWa741oZ3e60WoLZdcRXImjJJeoWuXB6Ng5doVX0j
SbN5aasO+neL9ein62+6pwwOC8QhQUpw+3FfeHpExKn7kRKqcyuzl8G4OYbOFPwY
bTNWVLR4N/dXSBekFpTWuQqwirhehcd81PTs/qr/RueJfz433V5tCJjIFv+6kih0
GjLi4VbzTZ49FLmxqHYpVzb29KQcl6+zVChVYyIx2b6rDZ0KDDm+g+1eTweHPBMN
/YgX1XVn00pPVCT9R08Vsmd1ybdDTVevQNqhZ4bSZB9B/Qv3K6vX4rmrsKnS4tTo
BVrTpTWLJwm9z78MhKcmQt3gAbtTsxmU8vCJ0ZmuVAZfRwBZN90AnEhNBcle00Uv
5yLAtz/sEgGMK6PHEBy1cKNMyYHv8/NYDZtayWB5LOou1PCEeKtVXWoj28BqTNFi
1CfoqtGcm47CozWEu134ZpRPSEIJMSXKrw2EXOEdx13DwtrR9N/wVeo/odH2z7G8
QIGP+rGfRsRyGCo6Q0vTy8+fq0pffshvqfNwboUz/2Y9rrpYbyi67EFYoc+tZQGF
v+GVMHdVVBMnFqa1dhUjfKbJ8nTvN1LBSRBKqqCFV9m9jDiuxg9AHC3TD7MCQVQC
Rtryw6rTSbwVkwmm6uEr+SfIm22FvEug8axcnld5kZwHg3HRKnQXsgypCa2Nyecj
G1f0tgM9Qzfv7Z4m7sIC8A4mAtt3OxJiJXj+4ley5NTkVfZKP5rGp6Md5tpuXRXT
Z04SNbmWRWUb+KBL2bmzwZW92ll5cIE/X5iRYU57EcUK9C+rQAEVRIKY0X9lFI9p
b/v02Qa52l3S3rAn0iJwhBRcuF8mippMwpPJRcWiExO9KZ6camC+88RSHBTPkvQf
EBX44y4EuDGfF0FqF6yGKcHDRa2fw0b/gxyxuIXRnMH6EpCB3/iThFbvO63+y38o
0Tn9oq9itZSHmP3ZAsircqQ7ImVO40TK4o5DhZbGX+VMoO5aVh8dMuW8QDJ/tcfN
jYr2OkWaGzsVbKX6E0vx29fE9BfJs0C4R070YdxtlcqxUWsHt7D3IV5s2AtZuf73
Toe5PP7MkdXOH7R4PdRbGhWj7Ac2aCOtYWygtPSfHN6Nks5fN7ppUFwouzbwHKDc
Beh9BcH07qEfOWNMCDk3+fJlIRat4k1wckVBVqSq30DuZRvLKiffZJ7OQ9nDVWG8
LHHIqO0p2n39sdhLqWR/3wLSSiGIDZ0C1hbrY7DBRl4f6s+6mnL1uanaAkLitwDu
pj3XOPfFtuf7mGVolZrkOCIWYEu2ES5S6dCz9YWK5ZxXENEfdYcdaa1103dkggHf
9OtViWy46F6Q+TZoZiljgphbcD1jELeE7bKmQMBYaqN4V3cxa0KHa6qHpYvBIN3t
kKmRaJbeXCK9XPPbbImXt9yw4+gTsIEwIcSvomomhojSBNokAPpcd19vcQ2YRbzk
bw2B2CR2RTLLbkCoKFYylufcT7VdDLgteOBsTnKXRFTYCuAE845Pj5Tnh6NPGuPZ
WDDAA//j4vCIzRWzi5sLj0IUTAyLvy3qdcLJnzI3ra/GlrY+8kViR+4Rw6cS5Rdi
4GgUs6tumD2YiYJzzhbbJl4BucZpzsjUyBgivtD6h74zjC9zJ7MRRgD2HaS74x00
FiPkj9uBj5czEvZGLYlzquCGK5IMrt3WqlS/oC9rkob7irOibkGL9W9dOYu8jsRd
bley7uvGdFzyh/mQtba6ADpC5sG7rNxt7erDULY5wvhaRUHkFDHX8r45hh/J2B1q
TbqKg3uV89OhKDiBZo86uvO0XinCvrjBIZ9JbgxTqtEm7P4BJOPfCg5Zhd1AntU5
bBqlfLDn5LnCMpCygoJt/kM5TzWBd3DUWsqK4IuKsHZ/9WVyxchWYHMav7KnHgT9
baOaR3sfqZ3FRSGC6ovJKXbmeQNdsrhTj9RPS1Z9LhCnk/lcyedGK69dIjEZ7NAL
R75C1ZIgtUVzeOM+YlkkW3cOYd98jnegwrRLUY8d0JT/w0MJ4ClUAmA3p92kd2lf
Cx4t4M6ZQBJPzGjwXdmaehipaIBJpxk6nf+ie5Hq2/1C7RvhIC8aBUMMfbmll+wF
DYi/9lN6BFuiAzA/6ze5Z+4wXq++vs/QJtmoNEQPWUh453flkO8KwlDfkj5wYwOD
rjo1KT8HOMIJURSe38R2xmJkpDTHH9R6tVSq4SGCe4/rUe41RIXmc5Ie7SdnGzfE
XU+Brk0MYZb1sJRZTg+WYiIRpB6VYZSXk3VzRKuKxycAL4elf2UY/eJ87O1HyzuQ
LFoeVo5rrSRxgGnMv/9spWXRCNzRLN5OAbFkt6yY8jcDuNYZ5n74WgF/XzVcK+9n
Z5WZiwQ7gZhESZSVdrO1KGPmQXrc3s/uG8LWc1MVoqYumbAQ6cMEPzFKwT6B6pR4
dWVUVS5jG0LWMEsi/JuBr6BUzA81gbC9+vZK/aSOoqPnHMq8eRGGaA3uDMfftVuu
EvdrP/J5jS5ZqRT0sggFam2dTTqIfpHdU9uOrekgQQ0L+fy6tAx1yPRyqdubrM7b
Qr5CJHIG9Qj8lRFzMGZhLnDKfFWS7wnIVmrSJV4/aabN9ri3vUU9uq8Wg+GPd12b
tGZ2f2QiTho26Tqk9kOLVmwqDomZIDJl8dD+yVETcJdaa/w6MfyVmkeZOXYTrKNm
pu/mMia8fvgQqpmgjrhWO3KgcHxdi9BVPvHKL/sXRPUJ+6Unebl7Xh3BD3VvgYcE
2N5QF1xbESy/uLKLTRjHJo4yjUkBQxoR6FpzF+pTcbOwHlNLv/frbNYZuBQJQjx7
3W1xIiNyR96B6EsN0TKfy1jvZqIf/uobsUR+FMveRDdVHOSO4Ku7g1l0LBPw3nqN
bGDQoR+J5B3TK7k378BC38OqMcA0fA2YpZZfhEtxbbz8SwQ1nVTCZnwK9KgNLaFN
TX0Upz0BhucytwwrWp9Zj89RKe6oKIrK5L48fUqqVu5zNwJjt/GhwearSR6aK96r
vb9wWCgLM+OdYGNMa/TDLHLoFYDjHTcOLICZwvcR/ovKK/C3xz2NpNrooD7NhlPg
7ueb+sFt9iSeKtOT3bhuF94fH0gLz30ShpHRstKt70q77rwajgB8XT5p0HcS5KZB
JraymnSLpB2f720ZxloBIjEtl7FpiIIXQnFdhtvN7Jt3nYpyeY73iQndbtQ55aQS
V9Hx4LrDCq/7EOrOpZueX8BqLQO6pW2i5pHS1aP1XiOvaAtUaSzuO4mEViobjkJ7
dquePALN7ZdZ4eh4+4lrStAiG93CZhS3dS9N2PVISZCUqs042L9tTT7b+Vs14P5H
J351F9OXv7pvzTZwTv6W869BbIoszdEI5HWonwaEWsNXjIsOR/ILQNyWvqrG0NCq
sO57IT3qTkZFSEmOwHf/Yn4bG2PoNDGIx+auiSWEuIYc+M7atMi1P+ZswaDPa2BG
pjR3ilN7NlcUWP4TtzEMkshi9zAZir5r4fi2sngbZ7ETmNDgYLylJs1qjnJJsoir
+kABDydWixob2a93vyjDQHiSw4HjBpuw9fUwQo0aKPFL68O1RBYvNipLZNIHvH2s
vMaM/PJwA2669dFqfUNEejs42ZxxVQpQf6NT6vhUUij72E8yixEPhuJiQF7gFVzf
IN3NgHeyBZawqcmkzWhRhFwo9WaQbTP9lTp5DbdVbNCRqtdtM6pa+CdV6+AJxS58
tR3W3tIUy1IM5XU2Qyz2L2KnLakAHm/TFmkjHVvYWY8ZbZgQH47aVRhS2ZtjwKSq
hECGH8d/UB8DHoD7DuOQFqAArEd4QXifrcJhBkel8y5lh8P+ZnRTpzpTZcirHrVA
6QU/osG3rhbfQe6V9RziaXo2xwDDNNzNAU41rJz99mOJoC3bo4cmbvy058+8kh+4
EbMcv3Bpiqk1V849rdtA5iX2pvkwvMdJVdNHibNR3wDj/QtYoGL/FbBqafZ/KtW6
A+PofSCs4/Wl/LXwxtDKuwiDqqmEGeH2PDV7Jc8NvFCT/kzlUz3q8ORoNCkry6Hu
eJF1h3lUIuFQWc9LdI8XCxk6cb3mtUkbxCHJCzk9oQNkkVKJMPlWHAipZZlrHoz4
cAWxPV52dnh8dghGNp2jKHVBcbBrP9uj8iC9tGkfWkmM4Nh4g7eNsv1PQCoL6akR
C5O4VduLFP9NQlXQQ5aEXH5akUEsfsQXOqKEgnXmNNbQUH7RMo8tDcgDtelhcxxb
vr9bpzezejIHD34sYiCMSsh76Rlv5ATDoNf5smvmLgZwd5dWva7+35HjyZK9DxB9
rC6R2LAzxt0+Duo1KImwebWERX8gHZW6xIxY2EHKWJpTuPK0HcsWUiYUCM577JbD
B2Nw/C2rHKELc6aX0PuBjBFKdf7zP2mBukdoU72eb/y9DOf0srhHcF5RIQmzQ1uj
EIZFtSS2CcqMfvAL2rnvgrcFFoXSvIV0XFwrqcvb8xtRGtKGIca/cfNSmUf5qpr2
iTdLirbdinZU/oJrfEvEwJeZ4ECSHdbZh3wjvTvh35TjgOxg7jqYfZDdK1FWv9xN
6WmP6nCmdabLBLdcbGpoeve/xIEftLbnil5aBKBknOAll3Sjmu/xO8zQsY2P/Z8p
/dZcIT3O9s7pzw+OTi9LFO1ugwP+E1lbeynKf6F99+kp/lmbcifhNHrTahjKQ7zW
vu32h9dwat4CZXXM1TfEvVeXPxV4JHnuQbzvxNd0EGR9CZ43uuxeoNH+WYFez3Xx
hRvdPVvrdbqfMypFnREvxzjwWd/BCxeSkcxZ3o38PE6xierFjg0iDI7o+3/3YGYN
yU9g8iCpkOQ9AYcUN06fAEleZeVwVcb/xmC/z4mOFta2j98glH2msIPELs9QSk3/
pE1+MGXe23PyUX1Nj2mQ90/kjz1tg0DVA9QHEcWGAd1wZcv9M23168F9GbR9TOSf
RYbe+FnFbOlacN1S8KtAmP4EUS095KX2EWRg+L6WMZc75fMrDRoko5woY4BVO5Bl
cyGcF/SYmSqEbIPxhjEJgyR2sadbbbmSios+rO5GPhfohbkfrK7xhsEZtHjjzE2F
1C9s3IqjvyRbd+hoXqM1Imkg4eW/Yhjphza829onOo25Gl+TBLG5SjxgWxCLTuNm
9C1DNinjGFCe4qyskxKlnbGqZhnCyUxbKumDzX15KFTvfIjfHQB5xMjj3PC/iFSA
pZEdkVoZXIj40sDAd4PQ7xlERzpJZn4TxlQbYTRk5K/kE1SvNAaGmvCxmn+MJ5G8
9eEDdSdh8l0MntEctzS/eIQ4WMGXHXOTrjCkT7Ibb6Jk5eMvZn0lSRk1xwG6nIE6
6H614TWviXvnd9lIrjYHXgkyPG4Nc2+t+08oMuZ1dloRQvX3C97xi1YTAATVRheN
CwqG/V/2hSqMTG8kLfKc5/QNSMOZTyP3dLb96fYPF0NpKzvdWzSDgpzC5dxeyMhP
GSjjaq9UMmct9tubY6PKgtu/gy+6mKIGVNKj4LCmuZTE3PsqkDERTtNhUSN5neOd
0+w1sKNJCzFZTn3bArV5CvfvgMJ3fzkTOJCOunKcKS3mnflPAz9X4aH+5ZYv7Kr/
0sqP3XqUlALgfQhpCBPrprUZepK+m7IuezIoVNaJGM46qbxRYXxPPGOB6FgFBW6H
Zp7/rLwRS7swiyqJnR0e7XDkQVZWnF3XskynnMLJlJ9TO/bky7rZECX7PXOB+Ogf
MN1YSRCNhpdaoZaYFxn45ylDbwyDDlD8FG1unCQ6DP2A4oKa2WjOIUsEYRLh9Euz
pCutgOWWm4PEhjmbnmmci1ZYaC8Iq91eMqXkQ8EFgRVmsx9fZ9V+NAkLjFqT7Tw4
2C98Ky4UeKGjHR13VgT/3jf1+A69lVWS/C2WQZFLmnjQEc9VPjSB5SHjDuRISyp7
THw+r0PtrH5BN+F2CLJXlvVg2Wv82LYTEf6Qw0KxOHBq6/5HartLgmmt0FDQa8Yn
RcfqSE+afKeXTco7d1OCRQ6+1m7PkOHUjwyWtvQhAOpaTTA8rYjr2SCGet36tscH
QjBBLBun+r2E/ka2DKDSn4DKEPS28oypp1t+IDhInOVj5ArfVIgXn4fKPWxQgEdE
gtyqh0AGU5zrsfgseS7WA2FmrwUsdCoBFOBOPnzdyD9AJ2LVq8Mk9Iy5d3E09LNl
r/97x2bPp1jFR/ZgQBAFZAnWuHnYfk7r2vW3TY/FJ7dRhlHJzko+uAQNVGcc5H+D
2HGItrPfKi0ciaDjRxobQ2iJ/EdJVyLh1TgQD56ZGnz7G6wtS4fOEFfy/Mjgh8nw
aUcNNm3hzpiMoVyMislByMQ6E3juGEtb0LnCnbARxlHIU3CY73RutqKvOV1Ln/g0
V5ip1kBgIeu1GJ0yuKzKBGSSDOECT6+B90iN/yy+pPabfzAHfyUEgug/USkMacHI
ItIWuF9pfjwhWttLnPXttfEGZqfCiFWt1WDukXmeMWHXgSFq9UTKilgu23j2f8g7
ieziwPJrnurhqeQw3P1DooUh+Y6BDLpNwvhS1hnuuvgys7R397S0Xz7sb3WpxTXB
V7ExhU5KgPeyS/WcFz93NkTTCFsp24JCCQct3hH+P3/O7fJ+jm4gPnpoC1S64jsi
rY+IwmYiKZcT0/JGcZYhESAUz00k9PVvAZ8oBYzJzab6ccNz5pDB9DoeKKnkIyNI
+DwJcrRPfoyt8ymTZ3IfVqPrN6y33ZEl1HMKGKzo/TltFNadR7R2oKzc87neQxFq
SNUrHA0WnAjph8Lit6h1ZcGCFEI9T3PIUWU+iSgVg3JKXwPO2gxXHeK5B/JoQu3W
9DRW8d1EOzQmTEF3XFJ9crWSkkClDxCvswKwzhWVtcSpuoaw6vshcCP1x+vI5o2W
CY9v8ak/DXzLXW4diH2nsYRp4XngUX2j2qzhz5vfcwdBsmdXFlc0e1GPVlFa4tG+
OIUPHRK4N2wkpYKZJBmdKPLUJtHVLrewGTa0bp1D2eDynz7FiRnzwJmI9helVonv
iVPxjtdqkg0iapM+TWTEec3ViH+VyIh+2fz8xnCqVPgWEtsaxS1uz689pYV+ZByo
xByzC+aZlm/4W5s1uGodBEQ4KnrtW1dyYlDCXv85+EDX6UIfhB5VZBS6fvDfTN+t
wxV2jNgkZudHjsgnHIDaT/27MpU5TMyKcp+LtAUByUUtTFLveXeidV8CC17lk9Ay
MetkEFjcSSZHVtQ7L3XJWkzzrBMG9H4eDlHuY0w8C+s5zZojS2qymy8Uf/NJm4Ia
sP3DPRr12ujEfqyHGEH3IIyme8zLO/py7myiHUo/4EC9hguvDCPMDWY4OYD/1fKE
SFYZPWjzjGLPBWc2armDA+8DU4Y67AfPLiQW1asykRgBB8TMXA/JkxOGqa8YD5pI
jjwIY9NpzSqpdHz9yD+8sGyFh3rzqm9k2KTOxyg0Fntu/eDDdQQHpXo65kvpo1rC
VHIEISNSOtoBbqgbAS+xXVf9/UNVVRNVQ4PwsbZC3g6Fijll76YgbbRo/zNpSvBl
PpekqNJokJshn7PL0MItldIY6FIREK5dRBvjrraGZSgPkiLwI6M5WjVcXeRDCcus
zylCxRoRxrlgZ1sp7FZ1MiZ/LjppXFIwqXZ88wgCwPLbshipnPFwWORFiK9n4YiM
Kcc0UCJ6YCWyfQSK1OZNgs/UoSU0ocq5QWLsmQdKACGz6MEyD3YjPPC+saSSBEAS
pzt/z+ActOeOk6NbYYzPyEOrCiFBMYp1uxiQeZMOZ6gQpd33xudr+UJRQS4cdtfR
n+YJwF4R2PC89n1EMZZlRpFzMLOC8AyUy3loX7HZx5d25GT6ABWlU3WtpX/2riEK
qwYXJ85w/kcMoPc6cE+3gqJMLs97ZBpwnwq7/UgVHL4bSvBZ8U51PBNw6utVLR8x
gYtFzv5RfHEOEdIZ1yk+enFzUYwDbVFkRT/njWmCWYYRjWR78ah9G1lKQS+r1T/T
RgsvIaF+4x5tTwW0cwGRso3BBLznmn6BjZEXlpsY0L5ggsVac9exPcq9zYMl/DyW
lXqB6JaIVBwoKM6vMTrqi6nlXvmj2ACH8V8NUJ4kyUvbe91k6Cs8BcyWRmcegYca
Y+UaAcIskWkiQGIEYU4QoVMSaNMmDlSAwHylZ2+xLpG3HXNMwNfd8BAX2ZyowB0O
87TnYA4dgLrT31CTtv1/NZIm3CzbU/Wq38XOiYJu8B3GH2MchBdAZ7smE/PHUHOL
rPdTYEwzrfFv6f5o+GjU1HlBesf9ftGQH6sq8zsmWYj8lmPNEflPw4zZEK1X0YCf
1te+u2bIMLKFR88JFf1G1Ms+5+/FNt2WvjiJzxuaJeq0cfkAZByzx1PCrJkdz2BH
6G4Du5GV2f1t3oQpKtztAExltbWha5wuAGZE/n6W0rqwS1VhkD4AP2z5Y2EZXQDg
5uXv6VLclITsOCdb0gZmYi9QcRrodjugRdadAid5B8Ems6lyPrMugOKAr8HwA5ML
dya/wd2fB/fyw343685uSYqHPPCri0f7t3CBZYZHtB01JXQHiwC7TOdGZlMDIw2G
pF+KfOZY3zVU1eNvrMbRptKBB9vuU/82dkoPGirzaac/XCJk39vlyFd8lLi8SHdj
h4XBpNYUw5VrP7RD0ed+ouVBUJ5FWHCWqQnaZKOE+D1xy/iZ1L58EHtsEKc4bb8n
qgeAX0KavuHiuEMLgIBUygyxjyP/WVG0ALIxSR5BdFkSzzMjzTjwgUHBrC3G7UwI
v9R/438gciiIWh9QZL02xiBhIvyaeW9C06mfmLa0MrWp61u2wYUwX906v9WIDQ3T
Tdwv4I5GxK7ylZHdacmyBCG+nMpmF+kqpNxPws6ka89XWzjhm0qGG60btsGOXwSh
YLdl9qryu31PUWoevUu/3sHqPG8qnxGfmsw3N3FCgFaUysiySDFkh12TV1BROwPJ
/9qV/vE+sjwEnOHK54KLTCMZc5C7glhWm6i4pvYh4JdvXJWjZ8pQQiLMgmW+oz+J
sxyEoLzA8xk7fKxNtufqxw5upBnOrUc2OUrFngD5heGWcOz+501124jrk/Gl5csl
jaJo4ULRk/J0Cjooy3MbWzwewPthHF7Id7WFUGDKEbAx1OgeRXLWV0nDuKMHKPhF
+UowkQeRroA2r2y1LKjUbIxcQI4IL3HTe0WD6o5Z6fPsjQHsI9nUcfl0+KcuSvSW
JGRqMKr9wYeXQCwZXqw3fchKvj5NcdjnSZd1zYJmRaM3wh2gK6NuhhIm69JuaieT
Sq92XqAeGPFJgzYxSz7+nlluv00dpyQVgemM8XXb8z53iGshQpU5lV0wzm52mltb
O4qxy7PAwBFvJ8TO6rixr0FGuC0+Y6001c+t0E9GWxI0QU95X8dRIM2lQSPjKOPO
+p8vptCiRmyWsUoMeAEhBvM0UybVyBC3wV7yxeAc/UVfmPazG57/acpdWsK2oYq3
Sb8pMFqYaycpSg3NXix2AlfpgacNJRv/TKBDE7ZtrIVC77RSUME50B7MB9A3ksLP
AFj1X3dA90X2Mo5g3+7JfITADYcVda1XvmuXED/3Bwk7b39fr/Y5M4V0SwbpsFeS
hgUN6wwv2wVjJMejFEppwIdP5bnU+q3JnieSodv3wZWwXDH5K6G1T2DsiEOPY1+V
pgdynWs1PoJOoyeUa3/FB1ZeUIDM5ro9DPaUU2BGpqp/f7oasKgaB28ZvmGko0MB
WIp8QXxEY6rCktqjAT0seJJIy3XMm1JlZ1/apHAA2jboZqigpUmvgdmRBhNzA9Oy
Yr0o9TODcGldb7S0HCsgOXBRYbtnrDgVPrE15GsHNQpfhcZWemuWASD+DwqnxCnN
A4Aav0+DRdw+WOPcqU/BmQmba1JnbVuZ1YJdxmo9196iBPyLbsHKaS8XcM6xLQsZ
mfwAXt0jQlbUAcjvqzKDynBECwd9aNBqtMwUKMRHU4sd1jwegALLljwytJrtvcuy
6H3Gg2MJ7tVlgJ9yxyKd5cypINPZifBuYqFw7MdIfv6Kpj+vg4xtVh3uxMvtubRm
iPw0fIIlD5zitqAFhdrK32V7u/E5tb60gNWeElLLOoCTszXcWQkk39QT9cfxQO4f
YLAtQxyF5KZSeV5cNcqX4bzsa7TXTl47tlyT2yLOmLOvfUTJdPlUZWxi1lzxdeOb
IQfJDY09VTM85YtcC1heyKRtjzSd45GvH8L+BrGaudzdZcBckWp3KCS2BMv0HDqB
V9K7Lgk93up+zJXfCCLW6Dy6SKn7LGibtdSs4nOnAQp1wLvpbH9jP/Me6xBbdXsx
ESYix33Pz3BSNFkxFZTlkIIzI0wSy71RXQDn1PC+C6TjcMcwFCZDdqSsb/qNJ5ED
kTULKFMvpRzGOaQJ+U8VfTI1hbhK/GDGTVKFPzTYNlpVlg48fLNkQU7ZthLLAE2X
iwPvqYv3ugNlruTxIik0HhKQ/KDUyKdLVZiw64AXUnmuMjRmgRC7uDm0WLGSr/E3
GuBDl7oZv087oPBW+7XdrVpGErv+cnnDqjvBGcSWIE6H48kWtXfWSGcZSAIXPoKB
Gu6jyfrUj8coLKVU+2yWT3vh+ojWIDNabIyX7qFcED3FU28xtpB/TCP280sF6sk1
MqdGQQ/1pg9ruy/0bIthQRIK/V9+wXpKHvzn29PJzy1KTppiRpi5ruKYzY6J6q1/
Pbpc26jtM4bq20Tcynoi+M/n2uMRCjrubj81JqOhRNGzC2LoRXxPkKsW0mhHTioW
5Fe1IUw2AkX7cUWxVINgYekS8wVEe9UMo4Gz7J9wbETl3iNPP7GcLOvF/6sh1KPN
koPiSdtcdJXoqYU09/3JBI8itarygN1AcccbVl416zVLFirzUTRZ68rUlfJicByy
WyHtuy7inLtwZvp126ZknDjp7TcxGykVIjEQtoc0C08LhJPZxiV552v4gUqOpoX/
1CFC2lasEPfsPYbe/8nqM9NP0qDbQ+8PC+fR1Kk+kKWqRgh5+D0kH2dRWDtKY4ib
a3rBtQrNbL9jFRncQj0gAby7txd+ARsGm22VSaHpnDY2ZhgjIAU2OgOj0+7+ojaq
fplrSCI4FdXVL/5x5IvJlb53ANnLl+RlRja9e8onSSHTQwVgvgKo6he/3xqJEchs
JttrULos6CJQjJ1BYjTQqtOwdIvQL/GSnBSERmHIu0t+VXrL+22f3YrhWQ9gyYxI
PMJXJzduD+PaKgU6MZwog7A96pPSCkW4Qi3DbOaORJqxW3itou0R3N3a9DLjze4E
esKataTuRn6WFWo9KlLx2urXQ3GiUVgbSnRZH4vEFnn94+NWS7AIFuzw2v+yfV99
1S+d8fBcJ+i9gOAB9I/bmIcXOjVr0iXJR7cUBLpRwHlOppj7WvIwRR4VE4o9vcrR
T2o+0tWRcxpOhcsXCXY8kpNVUK+JNnrHsKLQeFWLCYwLmhBR0yN0WtsSbbkjfal4
9/dhP6CUIwkIJd36oB/w1TYYxe4zeUKfW75dP/T5IebSLlyCkNpg3+v8vYUomyWl
eq1dKJnSU1eOHJURsZJVR/BWCIJO1iWHSNOQHca1j+yy8A8ByCcyoxikTy+cmLMD
0vrmo/TkljB360RpxEfKpYxYdi4AVJA/qWsE232EiBQJbEDwatPHFte65pzCPssB
c4tEIjp5Gq9yWfR1bGiO1tZLhUgKxIIu5oUtKjg8VA/JI1YBYQPNTWI6/i1QRPh8
rO9qTsi8c0J//Ca87sijSvmi9x1Qpc2bfgb18pzR7BTbCrhKJkd6TbV8TXXQsrEq
SawPia7I9doh2teI1fVGzgxOeNJ/HEu9zhJCgGwhanajixZDGdVWyfLCadfxRe3U
WWtnUyyQabwt5xzlVB0z9XbLox38LTVaKewjDOYMbyIBayKvQ1q4VDdEY4ohgzk4
gk6JJF12jPsI4KT8T8b+qCPV2haB76kz02EtM9NM+Tu+BEeFxiOvaqCiYZPuSdZk
7h8oQqBDLq5fICE/VNW2uGrnsAwQpe1tTDjkOlvV9+8zEKLFBV5BdOF8ZiLSS+Rj
lRg7PUrCXURbS2dJjavm+NAN/s9GHtysTB5iHVu0A5+e32ozUtVDNEUWzJEZ2YgX
oESVtYkiqfD0oCfsAebHNbcAcXRWfeXdKTzfvZtbuihAByYpEAPbWATpIQ5Y4KuM
J4YGxZ4HzJcQwY5cJsB745iVLs+ateRqob1bYCDqqYsNISzpJHjU7LH/2w4FjsY3
NahVmSIMrgouMTtq8twZLstisom6ZqV/da5pCOz2nH9upm7JZuJCWJMtRC9ifAst
au1AOxL2i2AA3TsoUuNUT313LXCvDo6id1VY4FcWgqjpQ76rbrlXI7TWywqkZxSu
vJiimUoWxf55ogARTHlR6HgKa4Q3yBCPN8/o+ZbkY8qOElUaY4k21vgK4PSAdFJb
qnrJ1ozGoDXjH5yE8ummOrASRWj8EqQp8PlGYgghmB3Q1GNOoAcysb1ozMRtsMdp
RMp83DQuX7/KFpnT0AnsI6AELGmyrntuH5AdO75jnHq+ImFAirwFWBEd5DO+6jSY
rNx6bduaNPZBFnDXzCoCBR7jMc58M6NsEzWmLDMk+I3r2mEIxiOBHNkztEvOXD6S
EmBp+psUnnWExak5/U3ItNTJLfC9DEgStKxpLTp/ueWFQw54UJnjS6ZZL5mBtiiu
NcIEksfQb7ZG9ZEWAK1YwOC1p9P4dwsIGZGMdbi/Zby0p4Xqxq4A4qzUUA4LV+AH
iDFPfioE2QFbNFt2++zmzWIEFCzWZIkUBrpBLWlDo9iJxHZijqNc/sX5UFrQhubH
ocYojmDrumzjy9Be9Ba1uth2D+QvJRwbhA9JSUmGGfwHTEJAmEdXuti1s60NRhQM
64gRpt4+YONp7Be4eekIz452HJ0Z/TLtBLoaMtGz3fMlY5AE2RPrzDPixxSFET9u
wFgQfyu3WfULqxayungNA+7Kc1A4aDAyg6pL9vgi8CnUnd5jcnhFZuSJXuT0Al6V
MOYpGUEaBxlwqblNiDj/0OweVr3K3i9I3Mjv4/Cwn5SGVOqFQs3sQiHWFtkcokiM
mIrD7CE49HAHPn+msiRNkbH/ER/ikLw+CsSCVz+hYixZ7m2xWWtuAwJEWlMAOuYZ
cWiXW95iLh2/Fe9+3whFkkbLx7dvVG0L+tmFJM0qu1QpMlcCeEjV4gGYwzN//twe
So4v7w6OehlWknAmwjjvRTbW3WoARuWF8poy9ydrPBB8BjuNIiM2LFsCUIFd58nM
6kGh0oe6OKdq1eGgnVqCc4VRVLmPlbxjmF7gCITrqB2+qTunssJrNRtEoceKWjcI
Loa/S+4R4BgAS4X3nmoYyC7K3MLjfv15rjXRttUkj1lV1CxkXIKkv+twywheE2wZ
aer2ZYTd2ECMfNmsylk/CvVf1MiFW/pjYt3Py0UHmXwebltocORLcsPzZRK70454
zuSvWuQa1opS9KdJdIx9R5EBSbhmzXv0D5FTvWrr12Whe9IMP7ave1JJCnBo7Kla
prbPRlVCpckdIgZ+rC2eOHwxvjs/kAX6aj4H5sd1C9YXfzRVf4nnUquOYuUCKdNw
ITWIoPnbQKzMXrPp7gVFRsyHDbzVTEkVw68+seUlxy7dalQ0KmL6FPyEPPbLiYm8
oYVqGjnnTiK2fA7gwLgOmCKET2cQIFUUAjH9TA1julqiR+olyQ4neoUd3qZjK5lv
jgMsNpYoWxJshKBijtu4kA6SWJWPFgWT/VyjKsx/ccq2C+f0/d8YzmZh1P/xLNxQ
yVPznvZz2hUuirogHJyXqu+IMdFnnMFrBpGqTWfTHBViL6FqKbBxtywKFrNt+3zp
GxZloESckJC2/sIkVu4dvD7QYfvPhB/j6qSTJVx/rosMUR9FJtOSmDfkg+97wiWE
md4nn5ROFUmXIDNVwfkft4pkT/07yx9MMWqVSEDNtR7lT5/pko5YfW2mQX6yIWy0
hJ8i+yanbwFx7uhLQdG3i1qlw7xyTAkfFpDRCxyC6BM/n1rsRTCksjStRNOo9K5t
znLVzQc8MkGG+JhzShZmd3acFUEtDHFmQOwvUHBp58UDlP3WyT7D11By3m9vNqLu
q2CjXa/9gbnff83x4xPWHvXD+9HNwLRmMp5yxQthyD/NpzaqOhEg4liuO/sOby3U
f+XQn8N355PTbz2uSbNxUroPyIbalPpkPaRJAiWh92yFFO3jYMswlD6ah5e48phe
C8EWZvNuEVa3Db56/jX456q6FSbvRr0JUx5NB90DKSdE0J68Vuv9QWOj7+uJV6n4
xDSIf8CL8w82ffm/f5FSZuDQsraG44HdWE4IZf5iy3WQd7yITigd19tqdI2MCZJZ
nurhsTStKJV+h+gaxc7Ip43zs+jtex+N3QJbB30jQateJNd5NXU12671uupj866q
OaiJ9zisdjfiH/i7YANJKNOKIVitirG9MZHoGflbBDyqmLextrSAsFqzPjTUorua
g2DgZ3ND6DuRs7A05lGOqIiL3AMgVQhcbXdY/T1qhwgK0soJxsgn7bUbbnDEAJBt
OIiD8Tzf0yFEkjcUyEjtvw4nOGg8NV7bm+3+0+crHMiLRNuRe2vHbzuf73foI8zm
x4WFo6GH/iSSRzzhRKoz30F+YipBN2XSkH7Xu3OFZ6LMIVC/hy0M/qFpr4sWew0Z
dMUKWuXmroDvYcRNzpxGSQlEGw5YjoOsMc5NrC7CafkTBXePpRQhnpHQvDLJ1TFV
lccs1DyTCAsYXP0ngqWeIBiRFPshgLiBf5PnAZNVUcUi+3rnyNyWLNM06ZompSiW
EBWN1ouxsg5F6Aiam43YCk8J5Obz8r9FeC+2v4phzhFz5aiT9QY/qs5z8OYqc9I2
XfEG2InSLAgvjQxzltJoiH+uW9MRqxSx/EbQuiZeAjJ0KsYeja20i1rmEIIf9uL9
MqcNqnJits3TCeKGdWeLGPBDQkjJKGjHyGDF7bnm7iJXR56Fwayg3GgZJtSCFZlI
M1lQRd2Cq50f3VVVGAwJxziltuMMv6xsgFK30/akva7qIvJEoAI+HRiL9nEpwTZz
K7bp9rbpNzmh2FGpOCQYHLcdM/qCEB8Ww5Wch6mU9bPru4OBiMujWXnxy5snjcJv
T6JlAdXW7Gt3XDtogEi2vfHT2dpOG3vocJzGCu1xoUNwzIZR+8bhytPVv7ik6zim
7tVsXnapSkIHA8VMwv2cINaHKP9McC9LvXsEsBUF9KMuxnSFHrs6OOMgQTpI1Hz7
MWY82jv/CtDs5ExbRECL4QMOB6zsURrUok3YmIiWCsP4AH1vQuLkMRxqzN01CeHf
vinMQebySn1s/TS4m29uf35XlrgNQygkybDcYlJ7XNiYVDOLvA6vIjBMUxPmQs4I
SK7ZehwIRZHEOubwVq9TrNqnHu0B7xtZRJMPqxQPkDrZf9L7meYUCNnGlWIsFAQz
DANXJ32yKKO+jHcCBp/M9KTeeUTTBR/k5Ca/hicPV+WUTErPDTxnwlBT+/hN32bW
VaDUvkJLtaGtc0RPB2RUN/Jaw/PetyHOBVYz1tf1Oj+WGXOUShbKyhQJr3099O0o
VL44XR3UM2N5ZarSf82KbAyaknAxQeqQnMfxJAR0SfH7HzcoBanDV0ZwN+tlvzHj
DwrCG6dc1ITS0azFax2EiVw02/HRLB7V401JBE+Nmh+Ayvx6ieHGIQfxBGOa3sNT
89MsH+Nl/JcHv8aW110A+WPoI7NChiAbMoRxCITgdV2r5q6NOrvikTjH+3dyammG
kvk69yKmwvdJ2jMrzVB39bjkHaYkFpmRUMGWPBmckqBYq/hvAEpfYAA238w8O0w9
BhxUbArtetb8XR5xPDDgeOUxzxULK8ZIAc30kAJg+2h2gWUsIiYtkVqYjSldZx4Y
CVkq3t2Yq+teR140ec72EB+WRcx8bOynCGqIGSNibWx1h4XaqrMfJYq8nzS5iqet
NO7j1+5vgWb2TqGlAhjD6fv7FMKkG0k4wQkgjkCHJ6TJjGifp7uHoevmDbfOsOG1
C4+3+oLMVa1xevvYiV39bgw+M/2PiSWVpbVtPYA+KsUfp6PR3CazwHWwH15F7MIm
PIuRQIBig3lxGoFBwEmS3bdj+b3Xf6rOLDrKM3cdyb/DSdfw0stLJOzK4LpTeTg9
XFPH8KFE+JO6Nsp0lxTy2DvOMvoeLiIBYDjAnnftezY0ZltlO6j4oxuDKZi0SkM1
35yLfTZMvWKdMFzyODz5oZuCv11QFCe68DGbdnE9p3CXfyRmT9HINV0DprPxSic+
c9cjPok/M7Mu9VoyD4mp94HFhLr0VYF1G+kqQkmJQkWK8frLyhbihIJUd7rnCy0o
olQkZhm4ZMmLTzrt5KcYdG/hfGTa9M104Sqb0e4NRBquionfxPjICbnIIiXQXl3v
avuBpzBQvyUXwVdLDtlgCSCKYW8zA5dtE81mgMlvO9sVWYDnYAIvYU084FV0KQrP
MT5Zjt80LiW4mWvSkuSt/sCwDYrkze+EL9mBeJrCVfcE/q3W+6PFZNFv3CboEV2j
AeatGY9mqGWTXDku+jaopj5yqZajx/EWjDkpu2QobfvPGEUgOBBWo4RgzmuXp+zb
RUuzN/25jXQgQL5NOFCd0cPRd3VukEDvDCqTnORmdyc9jnfQxhmUnGZunftqfsId
H6jPGoRad72jw/XPAW1IxbKBbTbp3+ABEzMv6gUxfp2ZqpaDFlAF6cuViwalxoVa
lVEGGofyDQjFjlFRrnAHaoqGA+A0sESu2ikgJ2gbA93O5Fmma9e4gCNDbbU9ILZJ
rE1YhUDE9Is2aJUWGYhi7QT9weW45bEwCuWcAnE+OVivL6OsxtjhGDEAsuXDuc4u
7zRYbf3ImENc/jYPgI2XGrsvp0z75NTLniy/4Kr7L8xiB9dUumKXlNnkKu1G+z3q
3LuhwYoPO7oITAhaW7M/CkANjqbZ/vyvSFyV+bz+jZ2WwS79aizZdEfUwMVlO8Vy
G1HaLdWN/3QUG6Q2Wt5GLveLbn8A/6voSnfpZbsAluu6DDjNuuzlsOi2OkrHGWHG
WwLGFg/YcVjbi1l7jI+1x/u/XWlhyKdA5gcLZEOLH+W7y9avev9QJEBUVa9rSe7X
DmgPdwClb5dPMR2oBLqs+4TIsJr7TEhN7W5E6VmcFg1fpvGY11B395ZRyAVEfnUo
MAxxQw1rlb1p/yDr/YQwFQ==
//pragma protect end_data_block
//pragma protect digest_block
DIHDRppBkL6pN+wIByL/Y6mSbeU=
//pragma protect end_digest_block
//pragma protect end_protected
