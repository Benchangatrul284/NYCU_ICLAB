//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
JEUj4PjkGvtx11JzR5BlEMZ2Cf8DNZHvSg+92yuge2RzfDan1LJILzgc4EbUc6Ed
qbpzrWfrE8NXECLpjU84MNFYImhBMvIm0g/aHtn3HL63NUTGrMkqQS9AU6ZWYFUH
E9LaT2rGAMu0rEGErFu3rTg/+UBpl49gX2VhhwrivpodMLHmatvvMu0VIJW0bxfE
kBWSZjHNZWK+bkLfl6fXILs25u/Aj2e5SOmJ3MO9LeOKowuGVBkLkaCJ2l0Jfnpw
bcgoqERm47EbIdOzJntQJiLp8KuL02jOocA5efWFfO2xppz625XobiuTg0BnFufM
DTssMljvSUHDskB4SSLAqw==
//pragma protect end_key_block
//pragma protect digest_block
PXquX6MY77HrmaG0l8Vm17sPRio=
//pragma protect end_digest_block
//pragma protect data_block
56KtOG3s2Z7l+lXyCGBatHky+18ggEbLPLRap/YzfjNV/+LCyMp0Ge0HILoaVnSz
7bAR6LPEUJrlsMkEJn/IRKJS+wDqobCRuQLEQuRST0r4wPW1uPoHC4ok+BGyr6cJ
Cr1LjI1IYcEhNgB6hpVrIr8B9cotcNx8iQiTQn2IRozgt5K3uIcixgerbk7DEEY0
FuKQUtpulf1wZyHtS3Sgqo/ASTosb36DLmY+ueLDChD0OSigCXP9iy4k/7luMmVb
vKAY8VUgSh8dfy5g/vpH1L640s9LHYIhx+uoXKTBKeNVOJx+ax0r85YiA7Tfg5ws
WQp5jCGPhTIYCN8pDZLBKMas5w8cqgvAisjo5i1cbdmrF3mL1XU33Jpmgtu9EzOs
dz/MgfEAHICnEaQbvngaHA==
//pragma protect end_data_block
//pragma protect digest_block
YQlRbsXDMyQWUGO0n8d7MQsY+1w=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype.sv"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
chiRPM+tyiuMCz/7y4xkwFAvh/3rVn2Ilj/hawaviYmiCq3ziM+Im0Pmihvh2WCX
YfZm6SGiHcOrYlci+LcEtrhYDBdVi/Nk8mnyIhVWRQQmzcid8qArkTP9PPzzd+77
/HXEyquKEONNsEx4KZftnU2XOi7acR+KpUMYyQGNeam9jw+gp1XIbQ7XFgaGzxtM
D+ZmZJb/mLRO5zrufWRr0jxIkasyiBfMrI/WSR+9pCvdGrZoX9qStzyG/jPiy+lm
xYkVX3bqZFceHQ7YSgsA2OTyE16TlQVdBEsA3t9kJDHdQ4YxTAPprnEqDWYEAGzr
t817eud1q+TFbgGAQSffEw==
//pragma protect end_key_block
//pragma protect digest_block
xxMEwyK/7i/kQF1EdJMCqm0meCw=
//pragma protect end_digest_block
//pragma protect data_block
2tLk8XAaWxzARJgGRNREeFL7+SbVDQJiaz6gOkXEn7hDZD6JjFodUjBJw4E7hIFn
roqHgPxVZH3LfZYCXUXDlNp0bW8nJGGCX+Zk631KCJHGDJ9WYSneezFpREAiDJzc
6o+72KxsBr4sWB24bBhJ9SBZLi/l5A3mhZ0sMAqVkEqq6H0pv4lEnn4lp0yF8rft
BUbhe5FVffWkC9ec5WzA9ooZGjrM/YG4s1gOB2tmaL4hcpUxB0nSD/K7lq8aaWz/
R+KWR9b5NarZV45bHAs9cX7C2EMLofrKPtJdDbrs0P2UTn09k2NUnx+K7xoR02mk
7YlBYlRbfT41eFRIT92kBCcTjNDwKYvKbl4Y8xVEMEhV8iQUDexUb36SRYRyVuaa
1rVqqvPifONtx6Y/6WCoEWUadkIz/Jjr7vQQJmlohTuxM231MQUc/xR0SLR9X0Pf
GCtHQoVDfcq9VkjPLlwdGcmQ36+nPuXHwnuW14zQP/TvJZ109K3fYdzfUX/q2l7K
bgGMjH92u9KYqAfH2sw45ZPW8wS3SAQq2hjSV35v9XTsnbyz8ym4GKsj1i/yR371
33YDRZzoc/G9ZEJ8ABLER94EvlOcIKz9zqKG3iwOk1ci37jVitEKH/q5sgA8olHk
xzep9nLbpa+jPPdgIvzh0kW1NKn2wsBc9sSg/xciJGmIhiAT5fO0NejHJXt7/HvB
3jW79FLgBBhGLbGWnaVrOOXQCo9GoGdRXA/0XiLfBozB5fDAK02PaPAp4n1BhmzC
iqdITMWKLaWch1PVovk8UlO7OcbIIyvrQakmZqDWKiN9Q0Fbnz1EfA1Aw1Zkspy4
Pg2qY+jx61TsPFVy5kW8yJT4voMUfaqIy5cK4xXsgow+vduGq5IMLGEsWQfULnDe
bGOxKcrfgX51gzBjyCsIQE+H8eHW5Qot1EUG4UIpmFzvDNY5chm9yk70x3eGho59
KM8u/qDhqudEdbV4QjWIzfWhWf/vVbaH7fAVwha+1DH7fdMHh89+JyXKgVSuM/1Y
LmwlICqoxAxFKBrgSlthM2vDAOv4U9ijTonb9fm40I0GkrghKkaUtUi6mO4M+bF9
SrXdGncJbHPft8DqKFCYB2OF3YH5jRxGNNVOqmPo0DP4BEFeQJ4X7K4fKkt4ALbQ
XRcneJAkdrNp540kIzYdfPvszkZIPIbCoqPVkA37+UVqXseUgusM14ngk+NPkmo7
WDFn0QmnKwQ/9LHkS59W68uVK9tOXQrfzJ6ZFDWNeqs22dQDHHO+QJLvsA+vUhiu
x9D12Dx3Z94TJGjvmRBJ9mkKONRdq0ZDczwKmP4myHxkzoxWLGXg0TRNBsDuwyL2
XOgkH4gsjV8DDaaIYWttBQtxHlk1rbrW05rG3SmLyaZ2ndD5Ul7ZM0vJc/X8IbDL
mpkmlfIwe6e8MIbdzgqf9KyLEn463sP++g2cnRz0DEfoSsk+QSBfujWxphq1DPlu
pPp6mOhhf5te7hltkSF+FmxWQAZdwS58npVvdDdlAzZrQFkZCuqTWvwfeb7oEt6K
EFZhaz2iJ9Vf8KuftT5kjQPrzan+cDb8XpgrSpMxPC/SOPNSVH8REluJ1lWrxe7O
9Qu358Vbc6iFku5JZbC81PVTsKTm8s+tFGavh5vCsTW99f8NYPC5AmcPGAWvA6T/
aF+F0u8xXp2iogPi+7kMN4t05swgjITSPvisEGlM8vLrrpe5rttP7Y2abfi4eNYG
o0//MUxzgfECaPYpGevNHJQPTZi2KMf5QGkf3Z8iav1PyK92teVFtVd3TELu1Xlm
7AIlsvaLVKy+Q8tjApaC+ewsHOsqFNrhnrFqyaOkh9DfrmzkBUqdnL7p9pTe5vRz
j3h/mXtHNXN/IJ06J5E5yjxJ+r7v3wkQAc9DUyUoNkH2i5Zs6NnWf4Xj4Sm1Fb/i
0n6jIMq4SkRLl3Y0ZwRCCsGahUFtRa4EybZgvmL5McbNF1AQCwpO9vtMV1w3FTeG
my6i80Lh0r8OpP+c9dI+Fo9jvhTGpeUWvGXl89lp8rpmGhkZx32bGbJKkAI/BKDy
7k5/RQ8bTb/vZcjSwDN9M5ZYRn1v0MXIYH3Mrqbeb1ufcTINQE+hSsr2jeW1X7T6
h4uSwZATRQAsoSm2e+bZA1/XCPtUes0MavHehU+x8KzUbyPPL8N+leFepDHawEMJ
Houyv7MeJ5aRp/F1GsZkJQqiAocAi3q8HZ1QxLG6vGCTe5Q4jW+NClG0P4f4wDkF
inloTw8rIim33G6Hcl8FAZ3QI6E4+BQaghVF4Wx907GziFeFQMwM4Hcv1B2Eorhx
enq1bIP9HVMpL12qCGMP/oT/wa26mGqVgm5DEubnHIZZe/MXjJPhFYJmQeOH3cqe
O900vGZ0aj65bLnczQC7JZtTm41Cf9kMjqNiWMzcKjJsshzFD6fvT1ncIJSSBPmU
FTxWhUoCZxh566dJN3M+J2vG1aDJEXdBMwPgvI/68781cXd9tR+3mDdncExo3egm
f7OI9b2J0XRndS3reM6awB8TzNiy+qs0KP0RqS0lGdZ1+O3CTYFmxv/ltAuhBcRQ
3465Z9G5Bw8r1V/3sYHs56IqtowVRU3W/ip2rcqo/Pov08AawnZvoXvLTBNZ8hMT
MnOP/RqH5yPWsULzSWv9BnU8Nfk1btBET8F51u1O3EEy/dPWAxn8guZVHzqP66SJ
gkVzw/Quiu4b6xEWHaoYWtuM+lFWF+/tLVxjnhff66YM1fTC4IdCOXbW0axMwT7y
9DVm8xZawaFyA1I3LL919ivU7ChvwfHB4rhwALG4O2r083FRuUKniNRNesyqHc4q
vMUJ7MoSiTrl58iCLPbAmh91n6Y7IOqRPVTUbUMB2V7MLoBhnzqoVWq6p+uHW7ND
/Sk6u/18dLV42/wdBZVHvangVUAXdvvHgePTOpt3hh2eonEOQA37o9JbXmHD6unj
8tADQZnwsHCT0lFNlahK1BOZQub0VeqhrAsvFWF/bMdwpTSMXxIQf8B3bEbSAUHx
YBl4oMsXN0FxjPLBtKp058ZBSnndME6OSrF1kZayv6L+GI3JLbFHAV4gFljd4Tc+
q39gcHch9QyDCUybwIvYSC/xPpbFGmlLc1faCTdocGIv3KmiFauh6kzt5s9xBOI7
vIBEv2Nvf20vjhI9rPULe65+yxTLcLrvPo6ImXh2Fmgsoesv/7X58hwPN6fL/7uj
U+FfW88VlYcQ7AFo709WiuYGWFmz1RRBt8ouiola9+Gh5jAa4ZQ2KBSX0r4r43Jv
hLIC/zDpzHLj3Pg8HadUuYnsPs1ovjxmT5r/Ne0Vzlaxnu75osUrATuEG3p9QqHv
SdTydGEJh68aJfHvpOYm0lcEOay9ED8pkfD7QkM0tcFbeF8+08rTXOf/MYjVi8YX
3NJ+yu0fWr004ms/0IFQFqXqTTJKbf7SlQr2U27xaHY/j6YopETWbf/d0XP6RAc4
1OmhUMkg0B4wV+x0KfxgEkwm6wc1O9egy7qf4O8yM6/vqYxKWAZUAsZhebBThUng
uHLaJqOvOrOp416q4dX82J19EQzE25OrRQbdgE25Cw8KkhwWC4jwslnKDSOUbZo5
2ODbyETglx5vHca94b6z5facqxvuIUneA5jxUH7KdTtiEKIb9rl+rw6UYfHUfsED
8d6GKfZvw036Bbirrkr3jP3QhGGXCj8XP0s2xwiYE91I/q8LsxcrjH9V4kl08nc7
9DWRaaoibW91VeqxS1hf2Hxnf7lP64ExkulJNatBDHNCV52lGgKvOduE9CW7MpqC
5nF21HTCkRYWvsqew96mW8U1VihJEu4ml6IXbXXVeo0DFc5MvZCVMfx8+U17zo56
JlDJly5xXdRig9PfH7qYYaqW/QFloBK5g26cb007mbC56/LkuwLYFJAmxg2GlBLI
P32zHpsnFpKBX1ubUR1EpuEFaPoCFu8b6KI/lHWEjaeMKX1EnwAoB1d/IemPDuWf
jh4kDTe0a/PCm879VNLjBVJBJl/Sg1nh45VSs5lyqu8Q0fLNKLxNo2zCQflz77L6
XDQw3hkGyejNoIr+qcmn9nY/GImvJ+Ck+eSRN5ZLx2AS0hUigMk9XeyDLfexBvic
2Wu+Agel9/uvMU/6wuPFFUiM50MDYo5QAAGN6j5+mjp689fVpHRrrZgMzPqTafBr
fATBqGZYmA2Tam/1sbGmwy3TtnCoSGrVHoW7iWLVp+2VIIZViR9HWwlMDJe7JWgU
gpnx+voZ5aE9bL7t8cSzJQ3WAbEM9n0mNiYvBAl9OKiqm8eEpHOOdV+jRQFESwWg
LRvHN5sBUjF1wVGRTqM5Es1yTPMyu17RIDaqQ/3KDdouMQoB1ypqZQXxr0kzKTFc
igbu6XY3mUeWBLTS/TvRIFku6wQ/8H2HGn1dX8tBx7UWbSTnB6vs69y7UDUGqpZi
nQXIsVIbvXxid3HLb5pNvLPMDokcN8Xlp1fdlulMBOutejTjqb3S8Swd92YKkpno
WSS0Qcm5J4DOcxXhubEd5QxO+yby0ek8Zs4jcAYWgZ5QNTChz8B2XhZsFq/vPoaT
S85g6JMwICv9f7Za6V3pmJfCjLVPU49sYM6iYHhsA3X87Ny90ACQQE2onpA9iuYv
Qy4VRhNdeZBHEub7MtGmVfqL16SYA1CIPRUpaEgydXnUwZrSYDoREAznxjtkNXBS
MO5lCiPbvLAOBLPa2zX2wB8Euwl/GgNkt0CbHIFuVefeAw/qWgif2ZK3+fAeIY2X
I+quPNn2VOLB6gss5dyINV/IjNOKyBBH0+UJnqPM/7340Di2859t8v8whURSZtXG
tnwyDFOQhvkH+ai9JxreC0F0y5D9VX5nT17IdR/QYJI5rpHZ2pJVNAsJtElvRg3w
mSquMx+GtA5dDZNcJbCmxhud9VTlkjFfidri/qXaP03cC0OXLfxDkXPRI1gwlXFi
B4ESmoPKlYGt0Z/vMupimkKNhbmLZL9n71yJKF9FYcNRp1ov2FwYhAOE5XDgNj6j
M9bE0wlqGrezpo4/uELy8ZNOYvnn5I4eWxhcWxq5B4HC/NNdDFjjIIzy7UH/GweH
uwJZuffxNsK3qulCqMKAYQl3WhSNkrh8eSQJsMtliJx89Ch3GCUgBtZkfcPYm9VB
kzxryeguDuz9Fpjtg3leqT4rrOgRuSgqXqgEzIRUFi1a5YJAj0j7JPRLW6/qzxYQ
yfrfpcBc++E2PFeaPFaoqX70k8Hk5E+vlR+y2cfq4M0ZjnH2QUyDYWfQAc0N5+a4
8XflcS0OxiOoZAjgrn46jfmFijiDRtKX20Ke8VsrYUKBCHBuPFGyf5k7eUpndx5g
WatEaGIi7AfAU7iMq5tXQnqDGhxZniqfHdkIpochTfR6t5tH9htrimbktpirBH/y
QB0dzRMQd+rThiulMFP+4C+LUct4NPDWr6AHMMgN8rhEK+GIYgAa94GJmpY84KC6
wucBWK7n9XocrWEvLPKJCplfy3w+7bxgP7gT6dISzJGoHSLVPrpeO/sGXA13D1kt
3PDngYCOH0pO5F/AsNelrxxlhUuhvkT2Y3rg3x1jKoMCkOXOprp7dQVlnjR3iUE+
eCLp12+Z93f4H9Yj+FjuaYGr0dhHxYiAjIb/3D31eMV0wsdYcSU/OEGdsmIJIsWb
0ndjr8tdTahf1t2mLJxXbmp0XDoMnDc6tMl4ut5aP/O92eFaTMmh9rxtNDZPqDy8
sIT6Bl7bWuO/K5bpqQQTgw/Nq9MnOvYOC0KVvELOgyT47MqWiYHVXZoLgMQBtmZ7
N/qhJcHtI1Ubs2Mkg1GTq6apLWzDzuUNa3YQD9S2oLhitZWTeO7W474N/Yq5Ap+0
zxpzkeE/Osx75ZAjPZjF8S0bRWE75AhsD7JOOJVd3k4KQA00QDxCfLLfPx6clMTP
C3XSW0G8MhRvmTZdlUvQo99tjoeYzk7ila9xpp2vVyzjZgJJKMdB2ye8Wl2UYfAc
qtYEGIj0qz5kgBhYy599ftiZ/Bx+NzVfMxzWSlr0IOtXnVMffUhnEQ91IR+AluvX
LejrCvfItmYpx5bvkntQgkukP153hiNBnvBtAGqbhe97QxMXboD5Crad9b6YcDgx
eWy1daNNS8GxjNzY/YMEGG+i+SL8PbGCmqMS62lgyTLYuDk1E306TnfiMiN8aw00
fsgZIRva5zO+Zrp+RxS+HVtTlXKbqOyqknYTld2x+C7sZC3MHEy4RT+t7uN0oY8u
dcmSkn6MdROBz1LFGrtCgRJOR5YqLVFznoVzrwla5hFxD7CYFoAqV7iadgbo8e9M
B6TG+avxDlqm+0qfnYAhb1RKqEMyVZ8cMkD8TKyHxcv0APesjpT6LCGdbmr7+Luo
UZd1WajB8udf4PMyd3qNUzdK3GbzxEMkLKQdB/XHKc/ZurKMBPCkh1SfN/Gfy41Q
vvK7WfHZO7PCMRGb2TPZI0JtVy3McG1S5ItbeZUKbbMGYlQ46SfuIL+5gpafpxQF
s2bXyKnMdQKN/nqweD2t8C3tE+wR+kRSTd9T0pwJiBjtei2y/W3cSqWYEHqCPGfu
BiVMgZu+mtYczli7KeRQjkvn46Kfx+/fza6mLHz2Y1d7TB3nlbx4+bUaTfwYTBDA
ZV4xrbVLncoTYw1CSjNpSp6vguEnrgaI+fgCRwiN3MmRNUry93Sk5lbAS8U34ibj
TujajM2mF4QG4DoXScDjXE/hPfEU4EtOpr4YodxolXLDYYJt5NkhtVYVwol7c/XQ
34+jN8nX1Cv33uDXpX+722CatqoAMT+k8tJ2wBKnldcLiJYz/IYaycBuXTURqII4
kOVEzpzj50bp9YIMrAJkoCyFpa/eemD+/BdhC4w8lg4nq97kLh+b1IhX3bwj9wEA
utSzkzPMX/kguDQldE9fyep2Aj0DndbA4Q26oxaE5E2l2wNzdsIAYl3azx7cNMSw
1a6lt1SCmstv24tSV0nHN8Fapj4LAEBeKiclQ5fmu46oDzwG/DVat60AAyqNG1NK
Rhx/OPpUsXFd+OQHSy86TvmGcx3ii70aWP8bzv+OLkBu8JNiAukG6QtWsnwgU+yT
CuOt30vvRZgGQVNi8KAq61HNPSNqY0H7NnLAU3NkDtKcJ2zVRO3wTM9EJZ+Setwh
UomtY1OJpaAT4z4k1ryYdjZvqFxJaQP7TNxtzG4+N+17JvV7o+NMCrF93p6GnNEx
Y+cYpXbeHZgYd2Zfrmys/hnjDLlrQlVGOEA0P28gZzgHa7wzhtFvNG6BaN4TLiYA
4yTfKhEQmql2L9JZSwG5GkbkYb0F86CG4hBZWstGsUrxXuZM0rlLOIpxn9CealuO
m718AI6KIwkgwTGW6+c+9aYvFKp/7nNAnETpyjHUrUsGo88nblf8pEVe7iIEFGHZ
bLLgm7PsNY10WLVM/0bWh3aJyYp86+a5sYJt1UcBqdMCxcCJ5vNpHhyqZe39VymV
VwT+tHjQY65Nh2QOHlJ4pQs9m/vrujbuTymmAD8vG8HiJquRLrO3jvUkmKVdLjjD
Rf1SAnmt7Qh/nLH8TI4jupLokeogS31JQMZ8MX8o/YA01z2waoxN0pOxLrWbbDcB
0a2aHqCYqE892JrK13/iHkjZoJFUyw53hYVqEIOTpf/G0i/M1/8iV2Hs/hwGY0DF
AQNktMLOiqwukbObSlcBF/7ry9YtRkdfra7RyiRsuNEXSoEKLk/Vamav9FriJSjZ
lKD+ZAq75IcCWnq4MZVqZxAomlEaf9AoMGg2rBvVyUGwi3wGQBY1DFcuHSsyIldo
LLZWzGY6ZNU2y/0T9TaJ9y4wrt4H0BpSyIHiwYyl9Muuf4rpPRN4d+80R0S0FQM5
fN4TJ6J+Gn3mDPGrm0JX1/YCBzst4jom+8RNWmERu2y1ge711lOo718wjZ9cVbL5
puW/+61JZQ9AjRGyGfXZPSsmPpMafksAkKiQK6dLi2wJ0Oaf2TmXVvlGBEyaTjg1
CeqSHJGIyNC8s59at3CAc7pFXqMT/eKKhi3w1cKZ25LdE2yMbSBGpC+HL5iu5R9b
QPqS9uOJhp1j8Lk+cIx42bDsfFn9QEh2lUxWLZGsPyDWjZkhWKcunyeARmPeB7W2
cRZNy/RtwjGID6aVdB3U1Y0eRyZ67TJ/ujPgMbJ/8wYTelZw7gHIZnr2ZATYc/km
NsBBB8YDG6CMPhiV6K1L3wuCbJc6EBJTF/eR3O7f4ljWUaQS6/aWXlLf3asO2qSc
zrYZ94ZUuYkDRIrC16KSrGMIic9MMCUXGP61c7A/tnrTVneZye+2pK0rl3U4IWtJ
KANLB4+k1LeiTP7qJ2Yxr2fHDdxL/19whOK82A7ZIeu1QM7HcJQcaP7JKiqYJrzd
TMwc8TknNFwsASkD+vpsR21V2m5WpXjOyJiX6XK2YWj2/qy4nc2HlRR3zMN6YvVV
9c43EZfWeVk1iKDo8zJngugk15Q0gsWgoogzWeYfu84f94qKlUCzCoW8eD17tmWG
SSETMLxZT+LtnFHl3Xf7hqBShy9sPQuAFEdEAenZjis84jJJgwrFjx7xsmfUuTmb
VYaQ+7ciAXEhB32UJLkTGlav9rTMstQQH9Ki6Fq/qpznqUQaal4hEiqKqubyJUwB
y1ALfgf03DnXAI0qTi+58eT9E9o2FzoS0xUirr8tR7l1frzoa0JgKo5LZpDmiRlt
oXZdXm6cqUcux2bY8WvE+CCGCAUuJT5XSmdzKt1orrJ82vVBViZczLF2QEhK8aJw
/aheBUcLdL5DRIqwEw3frHjluQP4pJ+IM4yoPa+LAG7wR3Pv/GizQiYwMSwOEN9r
mVncn1InaG9TS18JI2pXh8KCS1iKfIwbFqVqC4KP0KT3G6f14tHFL88CRB69Lgzg
Kfwg+SggabKlbq1sX0oCVA4P3eUCxIh04t4YQKRWp4MslYM36SngOepjs4ZvizP9
n9tiTleqSaMUmmoKELFHhsiU7md5XM2BE3N0dLTo9F+SAO4Gl4UYZ/Tm9tDeJSep
xejGnSTjOLr/9aP+HDPUB618E1vtLO0nnvMnD27eaPp5PXlUNFw0kmNycy6U/VQf
mn1JyC601Mk9AT42SaVmCd5tEf3hsP3w4K0EjpawloabzgOIt8fBbgOybVyDIOUj
2xV/uZJDBB/lr1JaD491FMO9EahH5Vq30hLqIGubfejKixeH5bsAYSmksf+ldD5c
jSxlAUpMVUiZhDxIn0KtsEtPNN4Ny3YQpWMSlryjiPerx8fIje7nYD+3rHn/Uc8O
Bh7jLFd2hSU2UxAwKP0m7ilXV9q4HTJLGZgtYx5H9lEHu4CLVevjnHn48/FcXsF7
5bPGY7idXUSTOvpjZUVkNuB7lFAyutYLQd8oqnlYZ6OCwCbmdqN6r4tC3pKfudmA
WUuFIC1yJ5H+aaAQMXblVyTPkHUuEeVVIghNwmQbcAjl2WI+GsTi4vIms6SMTwg5
9kchAFaTIJxQIGMwsdQfV7etroOI2l84ZaycmnHrFVnbtEoY4HStfCR8GTiPqsPS
nb5VNQz8J7AzJvtzq1V8j8flGL9bmhxLoABVoZmdRoGbu4Z20got2nF6SZYYk4kV
dXVcrpSQwHYAfdZKSMosdOWj5DBxRexp9oh8juUX7S1UVKT+df2Ck+5z9X2LVv9K
buMR1YCAjBdwHpr5WfTcBymZ4BjnHL2yTEtlXjdIrP9NBFmzlNWOS0UJFeoDRn86
g5Vx82CXlbohdhSoB8CUHpVYOAJT7uHdB8FQv+HSiz2SUSFYkz0rLq7cBsuPlpd1
sg+GwbfkjMGdYULFxmHMAKmG4iLgBXQ35w1c76Y6r7/wMPO2Jl0M3UvmltzarMJE
EM6Mvuundab8FaKsCzs8eBxZ//RNDJbeCC4LDKhOKFvLS0v+PIxpknIN179qKWX0
/qW0mDjkeUBlrFit33jLFDANbntDbB6uqbjDEiQhc4KNtHG0rSh14D5wqdfGaGFa
qdkS36vJNxTQdxrrVKVnx+AUzwXB+2xnJWaLGTg1SX98HNGd5C8XJoIWTbtwaBco
BRQ/QmGDUuuhOr6kxiImEIat4lx5eCD8BIM+PYKEmNBvhwnrwpSf9kgc/IN6IAga
CuEoi49K+COg5zI7AFCtPMqXQfG1cr6vJQKYkEZLSu2GSV/ZR3/35bL9PUe9cTv+
aZpdhGw4ujCeRpGqAzB0xvBABgE+ducvbp2OnRtqPPX0S8ooSHCDnvEZUdcoVK0j
fR8IqFy4Q6R/xMvch0BGSah+WIbEv89LTgoke6QAqxxNlhiiNVcWF0Q0smXJhGuz
ExIQIyF3qCwTahhyjqVdKS7jWCPNAxjsSHcwzH2efgYgqLMUgj1MnjKMQfE9sdbU
kCMiTHhcMNVRJOQxUhKazv0NoHRMdBEfMUEt/wqHgPsPeACaAIDJYAP+eVI8P3f8
s3wtiWUKxu0ZC88gPpKFZlicPczui7gxoPq/WeDCdby7BToRQ0yvSLpZ7EhhxIGG
GiCAQgb9QbSz8bE6s9jc7bdL8YfBpy8lhlXwpiuoEACQeBMP3qehqvKi7BHPOlEs
qZinkjKfhc/mDpz/jHuhu+WItMRa8lnOexFPm6qA1qoSBJk0AWlpMTC8P6bZ0SIc
KYCpwwtGOwpgnyHOpmGN1NDL6HxijGS4Z/lL7OXJ6QLCJNLJS5gaNIi6NYLmz1Gc
KgNQZWOQFrAlOkx324vOfn2Nwu2DvT52BhbQWmyjCyLjhTdJT3r8+bd0rXAV8I4j
PIgkubxGkcCjixd4BmRmiwEdb2AoefMzmuXUJJ/h7DHrqBtpaI3Upq9LfZDe0MHJ
h9qINWt55fwuyOjEUkmSNIrEOdzXeXl4bWXGpH49CxJwy4C3Q7F81gRNFYgxglvb
Ko2MtGnJB0CuFYh7ItSaQkzakDrzoQAwnLlY+gC2JR1m01a3Ckp86vYHluSS3TIw
3DiGsAiOdkIeW/NZxNEvgHe4P5e2155EhR5z1GVdB2+4R+QfNpX3ahNYz5ymxMbY
0R2/fQnvt210fEtAcZk+Y6/uJx5jK8TbkzBhhxAlQV4LqiEVRJnmGVsxn/fP2ERy
THVgA98pWhF8QsjlvjVDKB69nMR7Hi5a/YVn+HN1Xio87F4y9VC4h8RWhKv3UasS
mKmbEIcN0Ek+DJdl0t5E1F0nH/t9aNN9hLBn9gMc+/bpug1kbRPxFnXcMH6mUMgp
ttiBg1ysADASQ38joiVRPYK5K4JI9j07dShdym6Am4bSycEW7Il6K/kqfdtZhmDM
2mTQOgNAXMlALn78EdsmjebDCe8DZd4cxM/dpdVNP/7TcgnYQ0PQ//Ss0d5bTk8V
r7tnDLRVE/OLyaxeg5gAq1ToHxdmgCokn1ug0ItMX9TDahcJhFLh1sjYDYPF7h6T
msaxfTWruDJQwId+bQSU6bVExnQg67aMTL96NO21hXBvlXNTZatOKtJ1/OaDev7+
WNmjUWvlZl7lbcehMpDdtmKovn7N28vYlukL2nq9BjfB917uygMzRDHVyOefQnq6
pnQGsmYoN/qPvt2ogT1O7IrtvkDz6ClLuO7h4m1LE/duLYjq08rT/ODnZBacFO/O
NOSA1VDM8ib3oBqxH+PbFeR2zEKuiQcLKEmBZzgbSOjPAtzCvwZeK840+tL6BBFq
fEecVzz6vXTHNiJJQKwxwyw3CyKlQ9GRx5NvXUfWpww3eJfd/pMnDigqqOgOQ6MH
cRPOoNbaKaVuf/HaA0WKyfgxzv921xXlIKQ4FylRH8d5Lp+LacRf2W14NkWdp66T
sh3IYq52eUM1eFE3eerhgeDhjiMNTJWUkdajyBXe2/XpwT7XlDeCToXcc1FvokVk
X3UltJytbc5+oxCGNtBXm+bNoJ6fXTvsULBGCZu6cQgmRNcPDiKwQShtyIN1/UPB
DPB8gxJVNH6CDyojHgaNnYdh3yd61UchGK41zFxicfKjpgBh/h6Abb6zt7H2ku6R
DF1VL62q22u+bBTLtBQLnFhI/vm0CTNL1e9Fq95ZQeGcReAjRrBqDkYfegLIcwlf
cXHj/0syIm4KyRwJUU22oHcSL50q2Bx8k+0BAoViiNCzlJJOUFDzXCPK/GIGZBKX
TQg8MSFMrwG58JB5bPMvhe7PL0B/1bs5/kvNGf9dN5tAHzFzKOuIYv2T9j9Wo3fT
F2u9+isEYmfnCGMF5tGvFJdtBU4fL7k8ac7shLayb9PTgNmtvaH0n5G//EJCD9hG
SsVQsN2CbHw0Bhc8Z36JzRPNDmAiZMHJPASB+OzE8GCYLASNltIffmDzJjjs7SbE
GIrQE0bv+4/1D7MK5ltY/iYD06SU/tHSZmK13uHTvvwmzo0B0EMyNFP2gxWp5YvZ
1rz6aF72Trmx6cIeJ8FzMHnICfENvaf5nqg6SMGIWtyIVcTUpRh/02M+jgj7UEn4
3ORlDL1aLou+g8QobWa1hY2AzZtmM6deu6MlEH9RbMZyPLlu6sUaQIZZ531X/rcQ
CeUxMkCraMdPDhTUvyM0PEx8OVtaQvckBMXsdI+Bz47QvX5c4d1iGssRZIibUm9I
TwphgkHLN3mGpq+/DAhWGFza9rhjwfR9tVUALw4X/oKE7tenvOVwfBhy6KB5MGqC
CoC1GWAmcSIYW0okenSTKWvAEbpA9GeX+MXq83++3QMBdqp3+dzfFQRAblM2nHyo
fb+JFCwSflnspPipGXO9+N06keBeFkD+AmH27HFaOvZ7jrtozjsIJq/hUAEn5Qeo
Z7RCQxCmNG1ckhYLhafbogA83JTc56fGpUcQIWx58NQI2rpvMA97HfJAWDE1WVh3
Ju2aOPHXkTnmT2D8OzoVRNY3wIfcu45AGq9KsXAVXhjqN3uCdD075hWD3padM1Kb
z18T4E+7O2csSdILrqaYFotGkaKHVKKQ1M35wbxyI3/bWRhYyDUzQZvPZ39nHaoT
98SVzDP/Utrw1f5VV27Z3UAslr5Aybo5hYPvgF7klA3G1XowNwvp4kCMYIONkAEz
Gjq8MpPdROgZI5/iWkBAqhpxPMOoYo3JhxaG5K+M878P0o2OMOFDxINzAcw5IaDb
wWUYOLmyYbtJ/P7EY4oJ+DCnkuZQ/Z8WA1lfsIcwJZsXa1DJsX6Pz1Zw3lrsW1x0
X0aoFLi60AYL+ybHNyzHzzceAmfzrGd5nJ3612OIMXgpVaMdRA6i5Y4dMfm7DyrU
G5HG5ntdRONXlsRJRPmEN39jLgFFi2u3wLsyDZwq6PCBzOzMRySZ7O9flMfqMUwC
621m6u6MdAC9BK3rD4fttE+7NTjQqeWPHACZZoU9LQwong0SPHz8/E48rBIN1/rP
TyYEzQ2Y0xCMO4L5cqsWARCm8F3zNxBh3Zpv3uuN8037d/Bp7ND6pu8TAnjn4ray
DyjW07gN2qlem6PeEkWdwf3JHiobpkuo2ApQxZg23YWmxGzsFz+PlDpns06L1Uni
PBh8VBh//RNqLV2OXkTi4Wl4UO+C3Nc0iESr0qS6JvLudLdHhABfGnheR6Xq6keC
6m2SxYFdjTgXxj9M6eIMeSKO/I1EesuUcehfLyDA+PNWQHhsVPqHOBzmS9awWcsv
JcuAa3EfAoKEyM8qGXUQShYATt/SjjNYEIQNKWwTc3LfTXMMeIkIKrRkjh7j1UvB
kGwXLjgIu3eSOtE1DGJxaLc48lRXZa4Os6zobN+eBCxpNEOeHgmmTtpfDu3zjTcp
vyc6+ni87zSI1gmtVUNd7NoOStVKM3FnJyqt7Lq0jM+3klZsIF/BYEX8WcUtmxky
eB1qWPwmGRFzNI+JKDO78Bl/P6rOp1wE12cSQn9BtPEYyKZt9LiH/ylV735LsC4c
BzPlcgCgF32M2WFCWfV9aB1DnZHca4Xk3r3WVpztAqE0wTXrwhmG91L64AcFS1ZF
yldaMjNrtMLOz1rxMndDrO/GJCVnpLW4Jn/gkL30tvbvno2u53u3eArDIT2Vtuks
wNYKKEwYeleC/vVm1vHWe9C0UkwBifDhQ1omKfF12NU6vCVbXeGIAcZJsN1gtikN
vV2iEXfQhddBQ1kki87POSUVhMxVFp0QvJUNt1WKNFU751vxfPgQKjWkDILnJPzG
j2rsa80UdGO5q9yyuL/N1DpQ1tG+be5fEL+u9UUFtTPvYHILgwF+wVmIi/q4Y5pP
vHisoSs65hxn+rnExJxxF0/jCwkpnAdKJ3VCbCVePNefz/0OEy1a6KxIfWLXDGpO
faLGQQRXyzg8qbTphtNH+Cw8ufBip5jZnbSVVlTPUXcE/ct+R+QsqlOilqRUn/N8
VOf0wGLLWaPUW/8mqvkbw4PvPZ7gUuTLRbOO7i8vEq/p1RYTDLXNyBVqKFd+d4Io
1MuGcDqOoG56GMLMdgq6GDRlhPrOAXD0Y9ymo7g0Q2+kZIltn3GX8rrQfUUybI/0
R/UokCUtyBxaXfz5p36R8KBOBp+MfMh7wn8M+uZEP0X31qKQiJEwVXmeAkBNoq0M
TY0BCoOZ1zaiPtOzQL56MOtN6c/bYmnB2+OZ+8p98Yqg0CcW3rdW6apFqfxWqIsf
O5tSDLmXnG5wK1CZz18rIt4VXr2T+muC8dlTtWpDFrIExZaHC2JXP/0MvkVw8Q3W
8OEFsoko4O4FoEq5onAo1wkAKiH4qQNnNasxCcCmTXuXYCHGyxJLlZpflHipTsw6
MnHq/PXwn19wl9XW/KrnspEx1bK5ZlFiH7ghSOcljUd6AJBd6rXbwzI9BH3/pWKX
GsSBzwRksdT79wTFgXj76o6eRxiLk+XOwkyKDJxLTwweLJQdxMLkK39aiyYX+3oa
58UHi8pxGTZj3bfr9EhaA7QFmkbfzVg/iTFlcATe3d3FGoUni1HDYhA2JLUdSKsx
HCrLblRiYMZRaX6jmyoK0VxLMdU1x9ocnpQ+0eXH7pWhoHbinOwzWFdYtr9lMozr
YFW+CgEpvReYWxoxgYGW4SxMesu/3fC1ttQ3qplkpoJbk38Rwaz16+Wk7TGdQ6b7
T/6FdNW1CNwOslQahUi+O02hwfKclNiSKU1ullbdWBdo6NRpL/px0gZxb35u2F1O
z08Zrkj/IrdDmXQ+tkMt00fYuAlrkN3YN6yyjwt4FNTdBRQei6Qd+BBvBEz87Y2v
O9i2WQa55YYQBG0z1ijisfU1F36UsomMi3mDMEG7deYVOOruZz6LdP9ymO8EHdmH
EWL4hEoyU2vDnNWF6aoh71GHyWb//83QZdvf1xBKdPUMVDxXT5Ku7Dbi6Ki+isvK
3nXEvtqs5R92T3982QObBtHRUUu/Hfp6Pd8ZSiMB5obdnS3trRDHD4i4WgJJ0D8p
boVtU2GUj7egLudhaHokc2KqPRPxHsfLDzy2SFvypg8aLkdo6B1ReG2iPPuIP+tK
YVptB75w8uyIrDSvdPyTzLAahnNJE2FdZeSdRwmkqjAIb9wasJdnaUieqzeUPCEI
0p/X1bfroyHkq7W6vz2PE1/xGNCY3/U6sed7tGt4tg/WDx3KaclbpGS9uUh4J+Am
xAiLvTuEnxlZpZq8EnvhnL7LXS6od5Jw2J0L7q50XIQr6c2OuE81rxWZVUrPo0ai
cJwFQRO+ablhMWF6+zDnJAGZQq6ckM2P/lf3NeT/G9ObQX+zhtiHV4Ok4SX1sNhM
vJN9Iy545ZRBoO2g0nrgfWK6gt8wmgO0CQdMvQVnHHayhWrtc37XB/W/t5iVMEMy
DqOOfuX6qaOr7aMaULYA4W9YbckmCclgKqLDE808qgtQCbnGly7tP3QN54V4OqlX
+mu+KRLKgFpkKj5hRVRxu66V87+bvlthfmNCaDG4/FzNXzy6+q/wa/0zZa2iF7OX
lytZUMroGSoKTHMYAm/dBpFmXvS862mvi/3zBKVLn0xfGKoS9PFGGRHZETm+w6/Z
p0uBGks989OclOdUmC9WDsmnibbZf6lgPnQ6nSp5W70CkKajZEpTPfvTnkXKUSCQ
YaTiBKFW2A+ebQNfwJyxw4dgZZfQmL55n1LvNnnLZ2iaRxLyMOOt5E8cXr5d0GXI
jQMMPs7vTyWnavzhg+Lzx1yK4nwmpFgp9ZT/Kx+N9pk7TY+W6FjjWSEJ16BletOE
cbj9YoG9qcrVMyLry/+FTDBiKA5G2reXKlmhSsM7NX+EidPNis616eDlaCCAihHe
8j8uOlOyqZQD7CPn7Yfp7LSFnbWsJwebWeNQTkfjQocJkfhdnAi16AixGLI8CDx9
zP7ZYZxHfNmjwFN/ph18FQhE8jx+RPExM97+3Gm88gQaxrz5qVEDpp2yoGGYUEdi
6w5nYWBC1qCZCQ2FEYKR4hT2/6usglCNzyCMKQpBy3MJE35glZZacXHVydL8B04/
dJI8dsWG14lG1vPIAuRGPM12ZMooB3hLS5nirKAznLNTvsPrAMArLOD7PGPZt/1X
Gw3+q1xsV/a0gMt3b2SBhWqH0kQb1D19+YWEMx0FRZHKUiBBJXAKEqI8aA5aXFCr
IF1eyDfDHvRj0/oWGot9nC5GdhAvzNoyc19mD19sGF4rfou2fl3MLmej/wcI+H0O
tvdBy8myEeMMlLbuRcYRJujEvZGU5p6G2DZn+IVNqNpCuz6Oko2z6sEWgk4h2UqF
2fB7CwY2BAaXzJv6tNBkBi8BYrKWAtBTm08XCt+OkJEN2DFvbnFo0+CPUaLreB68
dLG3JMw9b7w0wZdv7HmtW5rOH189XT4ekjzwl8ZYtgruJw4KeWXAR3boKPhWOrt3
qpVbHQDKgQ3wM9HMqOk36OEluQsf1JwjIQZt2IRzEWyGK8h9UECvFypQa6c+eHwq
Xy+6ARH3fmerCxryD5ddXUwg9V9e6BVlB5qiB9Doz3sC1r4LFx9SDjHuK8OfmkM7
lJ5os8L+mOvZ8//WpiqcKNzKZglnlOTcOnrDsoKl0u29HsUrGZcWeTb56WW/5QNP
Lu+Sea0APvJ8eGYUgqIVaceER+fz2hiZmgb0okc3K39ExzR6h2Os5Sdkw+DTRLEF
IR++F27Tn892Pp61Me0Tnv1D4H95EHK8GqxciVHTEBieC7f/xwqaVcA21kW5V/0X
J1LHOssJglP5QpTm3li5dy0LPxQIiN6oRzf4BxbNxgpF9Gu6NtL2yt4Az8XvCm3M
Nhd/o9B6WwR0mZSSYPh9HN5e1IHnblu5BADKeXJ2yAKLdTeGO8E5nbU8/8CaxUz2
+cJh2ifKXkYmL+jfr1v4KF3A2cmWgjpnvrfFso/v6ppa4idrUIWTS9V+JgL9ANrj
YW11Te1etqTDBcJCo0fNP7+cL3U0hoc8G/yb5yVa783+nCcQPate4Ie1AfTCLSAE
9iUzWgtqcF6FykF3nTVcF+YzL+mg5iQxGGo1laYh+3Acw4GQHIwlDn/x98cpiyqA
jUzMK0QuvtVV/u/GY1xQ9mN9Af6p0M3AIuoVEu3zz3eA9Tpy1oadmT+Fb8ZYeu9r
LaBUH/0AQrmHwVzpaHNXRamHWzm2GPuvPPLYlmxGZ774SaG2ndPfT9sNqhHZeTtk
tBBOt57BSUzV7Bsk2Z2Zc7bqK/NHFNgu16+WfjiyvzogWCivaKKq68eoWbjlsi/M
sxf/UyOlHRP+zaXOpE9dlylZFZ1+IKLfxXbBg2rktFpzwpfY+UCetqBau5eoJPpV
ZGnL05iEQ+nCb+RNODfwz6SR82VLcMklX000CzMKa92+EqV03lyeRuPN60E9sUJx
u6OYswpnuX9neTzOwhN+0g6p4bZRFonnr8ojvCPCWAKv3uzKf3T4qPPvQfffgZeT
81oGEujY0Z/LQb+hWtsXpwsc7ft1q5sao+DTErD8E/ULZgWE1np6dtcQAbDQzfy7
bAYqqck84a3TwiDuxqss5NXD0PbXzKIv63ApbyXe7SO+bz3t1VkflhXnDkEkgV28
xOWz5ttzQ1xE5N/fFaih3DI+EkaXCg4PQmpvFglR2PFP84Ynt9pxKivXiLkJUTsm
ZVpy/2VLTLHVdbzruIeFOPw0KM5b1Y7AOI+7Bk5s5YlQOIO4F3agYUPbZ9TSxVOn
Mp+GJTirzHpyD1wlnswI5OVn/hjyHGd54t2ITWYpDC/hpuBXNATkLWQAEZhhoQ4p
2ekiBIgH9ldzacwZdawBPyinQwkAlT47TnbgglZHKc4W1ocPmwLDlEemOTE+Laxz
8G/Vpa78vojTri5ycj3cnJZu/cUfipFLGgUDdVYWk09+TLF61vezLY28/ww4NVcA
TRZ7F3mRNb8MS7sWghQxSSXEfon08so4WF85y56mQVdMy4oGPbfKYnE2XrZne02W
CgcJYAbnZz/ny0ZIO4YZpmIr0FmgqlrjXLWj/FFqIWcGyzmZ2WPqHpbw21kg9J4c
oizwKy2O4yJUG1KbaaIxIgFNznr/FrkfDnzndHEG7BeZ+VFCJXkpTpZmxQnXPWru
mPmaWPANQmmy+w4k8AiLv0BLsJMZmWN1owcjnsJ0DfGH7DaXy2+SqsfdQ9AGuDKz
3NLPV1ZA/YiY3gpC0H05Vzom2A0iaVrWWG1hPOk5ijqV+R9FCneJr9pHfDG99RvV
GCaRjNq97aZ5f0JcA3a3inug8EPxKkKkYgKn5A9INTtiVOMu4t4kpGDF21ge4uJM
z43CTJkzrFhN3YTWq5NM2Fh1OdxnqNQ/k5aWA16cBYu3jPuEalWFnn4djMG1MZXr
k++cs9KrYKjolVM1/HHrSBYt/Zn1Ujtq8qGDfnrsWcKtd1F4FUhIEpXfFDq+YOmb
JoaZbBfV1XkZbE7O0xh26WctQWLIthcV9FdwFVyGCDaSEG61eZ0lrkvHwfJp6QoX
1ADPv7Fjiox/0QWmn0Km8fxhtzKH7mRdECoPuwuaDMapJCZwjczxW+qvJFVGUK+i
7+TZDauc6WFmO6KxZnb9qSiPXQpCQit5saodCDYd1nnIY4K7hNyuxd1uTblB36ht
d6o4GPcqfaBbvEpUhTAVxtZzNXLdkDYfeSn30bMCIJUaDYKckUMSBVBSDy783ETz
JQhZUXqovF7crIVC3IHfN3Ry2EtxKbR12Wm1AhEGrhmYBFypLlEbHTLTLfUVfisp
8DJCjC6cmpvdUqJrXLf3gNGi3cpfQBbabgkUZNdg3Euc78lMzrak/OCYbZpanXOZ
1AbOQYQ8ilkSwCShlsVkBlixyGekdaGOtG2x6FSuOXJ/vygW9509q38Qpjo+g2lP
7dP54/khSpB4wZwcWLBM7iiBrp2NVep5ZPsge7kZsAu9xLJ4jI9MoJCgvmBUQgif
JwW59TKqKOQR3EAqXQUhH9NwgjSslW3+SmK3XeMjrDGhFZY+TwxHNm3TSuF/uU1i
8xJTeJ6qTavr4BV4W8iZO/oah6pmvat+5sdQbmgMgPa2D1rzZG53kAkrKPxx/hWm
g2n1NSX/oXRbxxpu/KDUY9bc6Suf7FabX5obijsfkWPcMYFDAwresCirzXlEoL+N
M4dChRUk/C4WCkxPR/+uEzwFiCNkeu5rz28i7By+Zlsc+UuMiT50hQavc0yNyJVT
lyw534I3fedz2IsmXoOv7uvfk1lyrTvYvdbfAzxCMRiVoNDgOh3MZ+g5YAYAxvd9
ohc/I7R3K8A9gEu3o4pyaOhz8BD3uPvTsHdSS/8Cti2eBIcVxIwwLcWCgu48n2Ag
OnQpQat3andFhkVl7+ATJ+lg18Z/2j//0zb/G6Xf/sTlmDDuHzuyvlyv2W8SUiNG
+xCGORS/HKx5wt2UPCqXxJRuo80XOcHLL0RZwcVCKx8P1OwENqvnqwhgo/+LPj93
NMK9NWJGQFgzJ1Flue2+RFefGB4HOh9Rv0GluqLm31OQU849ls477aretF0OBDYK
T9KDOH1QpqXO8N2SlwqX5+yTSOg+JaRp3z7z9+hNl6ctqwt0Z4JFFbF0+hZaF/3W
ss5crud9mtxSROmK2+2Qq4IeQwAMIWQ/0e/UQs1TgLrXtUbm9PvZ2QmngsXQOJhI
PI5LZb/DiO9doN4GD44x3rwp562Wm1nEILtKRNsWVRd2fnVgh3Epc/VESbvfAWwe
JE9SoWYrQ8fIYRI6PWzHQOH6xgw92f2XLS9ZRNsRoBkjc5wxBfpeJXbTQek6A51F
uba0lgCsjp/k7MBL1HJGYxkjFmWWi8vb+x7Wo62JmR2SWDhyWW9fs0/o5r2HFNn7
h3Rr19BhNExu0NeY6c0kCm3zKRWga0IiuPaRFcsup+MYaj05rT7ftX4jPCHgCQKF
MDdQ5ZHf7EHmq9+2S0jHCXgANxLA8JKu2iWH5rBax3ZldXzL6dK+c/2vn8iyfRu2
PcUWsotjuwhALl17rocvVap+B8A/Aeko5Lxd4HLRVqWZastwyHDbMGxZgLcvANbb
gdCtVHmPmL2tyPsXyBn4DZM0KvExmt/g0YOprXncSP1iaVC+SU7OP6ta2HDhhn2t
+aCIYRqtsJUarl6vSMSpP1c6aABOMleCHwm0EzxoWVT/FGks5fhagZnMt2GGlsE3
F8BYlLMRCTmH3O7Rv4y5hgYQhqNdqyEwcUYs/gsF5LPc7Hdr/AX1R7ZpKjct9f6i
2qU+IUinuHrWjl9QPH1j1xbWi5skCaCsoBKmGNdq3FBlancMSYMRzMi+GLt0CKT6
EYBYc8AqFzjJohRVW3JT4On9BhpJmc6wkZYQ0kg7ch/Qb2WqPYdyL4y8kLdcR9aV
eZC8uwhYI+4uKnJwM6x+Q4E55y0MIIFnhioIn1xsn1xMJ9xuBuz4+yzMkuP4kB+T
iQcLjPfCXtRvJmrxYvCjE5XRd2h+VcbOCeqjpm/IlH4g/gk7Rmt/O5v3bXL2N+eT
ws2+qZ8NpgdCc+HRTDnqy4oFRTpa6XAb4hLRVrrbG4qMgI9+kbp5xjxGDqJBitk0
bEsdMHS/fjRU4s3EN7z1VlyX7jOXOx1jEI/f/kEXBD4f745iEkgdTNx0ban6hi2K
y9o3GBEZQeRg1+rMJr2j2lupNw1X+lzSkHP8Tql5rGdjxAYZtykFcpv1M5XnLoxW
PJCV99lE9m9lgAKQb5WfQtXH7IS+ubFEg++VfKDyZTeVYBZklh5ytmQNB4RKh5OS
0VU4R2SvBu/zdOyUvwGRpJBOnDhzbt2SGqRRPnFlXyVF26HSBkcjyohMS4o9bgTX
Di4VRUkRryDd8y0qIjIham3hK34nkWVfFDKNv6bTqEKtN9kx9Y8dZbCaLsbixTD/
5Ak8e3CKbgjhcx4NzW6f1fdXoNiMYf9xaxpBQDilSQFS/turDjyhPxr20Fq0mdUx
PnMhzo7a42npG7u3XmnFD+RhiVBQIoWOiHUTJLUXjKzeeSsDJ6T391m++ctovek2
w9RtLnCoztP+eGy1dmObf3XtDxAH5sFHaigFRHW2lbLN7W4+TSNqzgVqwTjMoA1z
lwRm7a6z0ITE755zCwq4x83xJX7KGDmNmnEy3qGL4r+gukcs34H8fvLqx7y2TwQo
XC0ConbjkAtXsU8Lxt12jTYPYnFbIICwPVi3WrVGsDEKepegzQQLUdjiPQmHHdQJ
tQHqu9y1yM4E4eor9mc/PCyys6CY/670UcwWJGT+EwegGXMP0QSxAWRP4qasZnO9
JEYHYVOUFq55DBVgzH4Iv9utvT/qGhDazr1wa+9FmmyKfosc7xz0EO0NEGdzBmBa
JvhUyvCnPkrxKznzWYvjV61CCpbkGzfa29kjH2tQk31l1tAuFv4ol8DBivyGY3/0
UR1ZuDZbKDqYmzUqTP36H47ziIoIOafMSLZb4a0G3dKPDy6jv3NA1Cg4bEpUM7s/
rn2S75T9Jeb2G0AnrZEs1WGONzIoOuW4b9ksKqleL6GQCRFWs7XopNFsnsd8u+Y2
MukQ7rB+0Ntamy7Mjdvn9N0d15odwn+pebX+OzV0vRis2cS4doYTDp8and35zT7r
AlsgRXl0dZRCOYE5GaqfXObfs+EDOYqYNUKTo+I2HcEJQXTRvxi5SvoBHYtl+4h5
ZONYuZIFkCsZaFwyn45lTjvzBR1QRTSFlZ06qB+SX8rtHa3+NIz8dnY/F0H49DHS
Lvzw+IeJ//qmBJEQYs1CnXRvSd9XdxwAc90F0p5qANWhD881n5lX9pJWzcQ22AjD
IfYVNL+tjhocyJw7CmGqNQ4KoD9RUDfb54PCpOUVvu38jf2AYT2zK9sOUodN0JTw
diHrHODixbMbc1+GLN8+4JUW21z02JnYFA3K2zj4O1Bff1/Y95zpLeRPUsIVDes6
lPO3liDwNj9HdH6mPp/RNq0Hbjc8L/yCGuLNH7rYj34UsHpGyncRvM5DPPu/LMV9
aB9qOXvdyJvopbU68B7tDm0VbO7oRfFcwVq6ToAc3xnFSiRbij/JaoaL5BotNEfd
X5JLx29xHtV5qHlZVLqOsXW5M7K+31C+jKkhIlxg82Y7nlswszxHP8s2d/r2Wbas
xKw8MbZ85nRAQ9ZLxtevpZIt1CBcaLQwP9d4/OJVFd9KnNKHWMe0OeM3SvckVi3Y
m03cX7DHm2cttCLMkrfygmVzG9lu7dwwUxdnb2D1YXCt8zqfeBH/GSbXveucECke
qjzfWDMW6NgiINlyZ8WdYQHS3S2rENilAnMGjFmtGHU6RWUaWhD1JOmcdyeL7ChV
chObWVetq+ImSTklDHptrJmqg9xfBnAiRAj6iyR9fKdzvaWlwbcpk9QmIRZl1O/F
aKU30hhX0z2+OQT+Bs3NIwqMaU/w1tjXqUxBnOjMtL9URT8lkqPV5iwgQ5pXEfy1
vh7Wfkf2texMK23AyXkpcuq7zczxs/X0oNZRpl//iNqF0fCL4BvFdOky13IEn2j1
6FCbUVpfq7uSQlZLvyvKTTXjSYUvvq7kuJ2P0opC8ps1aKoNtN8B6a/F8K5O/cEq
hQm3XJ/EJTU6yBAcdKcuOCUrM7sCwHsTtjFjtCvHNyuj8vc50JJNsSAZNnNO25hV
mq9cKEkVWqXdhCVW4GNNUd4v8moOCjffzBg24vv+Kc93SVuIKQM9rGiryrLgWL8k
bXWzm2agymp71Snq/ebW1GOjvRxcFZMzpMVinTPundTVZtWAQSmNJE+nTcIXFwcp
r07OyDCP67lMUJtOO38INbDFAyt87x33+SsH73v5O0rG4CUOp92OQqxoIAZ0fGSa
7iiGBzayx1XAHrg76+DlhsuVnCGokhwY/Y7s8bQMuVnJwdqY5qzyok543tNG47EU
Zo78wnK7Aeh+wNKi+ursaP7hIiTEEGn9RVd9saLL/2IE+LAkhYtSxF2TugDtmfbh
n4Q3KzuJ0amu9WEGYUnsZmxUOVWuoWkyfU7oE+ABrfMPwbl9WgOO7NhUbt1HoHhn
X0N1bzDgRf0KiGeCxgkZNTvD0UA8WSb5mSjB0sOG+prdMebC86f3oynr23uHSAke
PCEqXKydns+iKBcT9qOTyyVTWCrOoyyQGOHSYA5hBsEycfOvWuE1XfhWrAeXvmfW
i12hIP7pgFQcSkXVa5TasGvHf+cFxoU6kJhgP+dsH/wZMfL+tT8WRiZA7XhjT3to
g38+h2M64bsGfuaRPs641nYjIGqZwDk5Sg/hHQaEy5tNhSg8ImSY7QedgoEe9JAk
Hs+Gj19BrOOfcvVBTrl/eioCwtGV/bHEA42OkEYQYOykdnxgaiADIL6KK7iYnPPz
YYZjD1jA8whVce3O0eBzOjIHdRzoaw8qsX1c976dA1XQCppomGAn5801wUXRKteU
dPxD4qIT37N+rTImjfi5j2tEAQkp1hPRBvE0mVHGUjPgDeir7ucPkT48ayA5yTko
m2YLOCFXFtCsFvauD8s0zTAxIHFcuV2/Wq0f55zKAg7LprJuKW7MnLEYE/UfXtzg
C5V0nWGQkz8/pHpdoBkLEvbc1fT05FGWaHEKbhIARuCE4tHPJ3c1liw2UoWRnSgF
xGbGDeqow2btc23GeOlqCQ9BO23HkIDcvfR+Yuc47iDVEYKD7R5sGrkaAKAl237t
ZfJNcj/sNnp+uVfavAbEuSUOEs+2k1nud7ylqllrB+6rgz6blujoUj/i1sm0MJjK
v0KokMtigtmOY3RQGkPwlimKLiK9WIiP62+lw6pizxCZggaSFbT+dvM73OLUE8PC
K5wGEHuuI9Hx0MARMII6PrSTQsgNEzMwpdwCefFyoQ8q79XzIQeQ+QtE6iwXOG4w
P0jP3CTfSXRMY2TcX0YAD4mrlE9unUpRLFUbOURPsQSx4Jr/W8lojRsg7l9MW2i7
3UOXakNUxhYDOw+GEYvzuUqFmC6biAilYv+JMq67kjK4O9EWmgkpCyswlI6P/Yal
C4iDtj6vfZiOPRwZTEPY37/LiQTn03yWznogD6rl/CxGdLlUaPcIGltRMx2BIXOU
j3MQYYdsZileYXyp5FGFswn7DwDq0Z9Lv9iGc5tSpmvPpLIjlX2+L+SZcpiVXKEm
IQ8/vgqw4Ro8RdKJeg34S/5A5PjnKwiYhnXzzFX4b1hENR7H88O9rfXH+yyO3p0O
Ed6fR34Lz1As6XOWCgeyofBZADZxHE1EgxZMXheuE3kEGxbc330OL8CvOLY+ReUU
iZUr8rQTE/0d4/soumCj57rQ9qpuEJZIVKdrAkXgdtvJRcVd97UP28F3Ji43uR+d
v7sDVwIlpFagR+R4WH1FGAYHE1mngvoYUHKcoO4Rn7qU81TMuiXb7OTZ/UcGtA96
9BwWD8fRjAZXR1005J6itW8aTvTVIpC+B/SO9Lmq1QGD6d3qRDiGX300hjfCcLms
pEHurDi5ci6M/Vv2LMdhluNG8ALMESkveddK+df7z1MzqcvSYVqMHXGs0eN0caGd
MKy3Ro1jzTdjRuu232i8wwnYTr9Lp+0XaVuSVcJRiWaTJ2NINfQu39HA2NEeRxEh
4AbtIASd7Z7huWmAX5Q9fYT2eMZ6WYv+TgN0ZC1MMlXLX0q56OV1yQu9RbfjVK6q
lPQgaLWyeFUesqguX6FyjxGXE/TQgFEYCYRRep/iZPrghFir9MZP90eSqQcKwkQG
GLRyGYZET59olC5hEFIKxK5id1uRq2pBEPYwYDHfTzpu9Qui7krYzWzxIYjcAess
/7gpE1g0Q9nG3fwBpigqjZqNNpLzf0a9JS3lhOeKzOyk357vYSrxYO3oMKDkCEIq
9jOEF77Z+Cn3SRpDTQoWdZLUg7l5R+Y+Vt0NSy7E2/qUhm8IuaH12kZ1yMxZ/cfp
DflvYfXfvdSCPXcuLBLXoHi4By4I+Wz8FKgefQO0KeinL0Hbr1iDWPW17NuT8/aW
yK+4qHeHYIpvYsF6HYhzs9RljaREAq4wWQ7Ob/AivP/MZkpvPPFcQqVjFhFlpzsC
mG//h2oJ6ppxvbpLGZ8dHUCcZrpbCGARVLfdBH9cphtX7bKwsmaKEn4zRCTbx4up
ukH7/zJZu6V89MP/6zeOjbWg23DyrCfWCCShm5OXeWqMjuSL56sJhOmiEwdu60uY
kSogegtarxx8acrqcvbssN5hCNwS5sPsIUKBfUxV0gToOZkudGi85gldEOHGgjOK
QXu1Qrj0gFweaJ30fht5BRyELui/UDjuyb2Z3Z8Ju6SSKHMXc6WkdXy3aWrOzEF3
crZs22WCGwKjyUEQ6N84KYlZDL0/U9YS7y4I8+H+bMrRvfFeVN0Wn56yGsj4U85E
TUqXylhu+BA8HhphNcgKD/JyaHj/SvZ8yF/FmOpz8mFghydkuVaHl8hg3tkF+ntZ
by9gr0W9QISQerB5P5EFjtH0tObzpMWT3Tp3ORSAiHQCWAaKGA34Xa5LXb0xnVdC
IdcaydndcmBsHPSdXfaZnr89RAMmVQOKvYtSRQam3Ymyhi4TcG5PwPzgMiK7cPGz
Gko+keF3J8/qwFusPwLPWMsM5dFlc+p6YOY1u/GWaip8jBaLai2F90r3VaAg6Hcp
Q5HwaQjNbHflC/ifUPu9zpFpi4jXH6hcm+L82zYvusaAK7M/4b1sgn1oEAxQdISj
WseOSAP+/LbUJR91QldJIxHH3nDDOyrq1+EozAeuGBHXh5Au/cdfkJ5ZOLZsw6Ju
Th2uQ7LoAbwtNbxvnvng/rvCn0zXYkho/IMWCfh9Mpm7DB7rDvxk5kfj+blnl/U8
aeYS4IQI7AUz052m+0n3IgNTM5+CuW4xbZ0UlNleZlk+o/Ne8ureeFKLGFxEwHzD
eKoKGTsDFLpSVNIXFFRq17WG4enV5IwRloVBY0g0qT8mDk9BNBbq3o2BxscDPM3i
rCn5PdQlTrFK/Av/OgkWK8a7Zhc18GtoQDD0/h5otBwn6Ux6PhZ4cLnPSzXTu+Wb
+pBDKPh68RUyxRdejeiywENgVc+1pwpPq3AKYBfpVDnqoaTU3wgnGiPTATIl226w
SOW8l3oh6jARQ7dsUFnXGekAIzJsT4yEIf60oYMsh3/D1hYyOnC/0G5GwB0ZF4bV
PEgq6ot9QRO0WPuBjfaiBkDKY6AfccuFxtoUYoWqK5kR0qkhmickA66MSKjrR2dP
GoOmWdCWUsTcRQM5FBODyMQSVnPdkD5jsHnVgGFZhL5NGDvPtlC2m4BuTx5EDHk1
qg6cDI0QXtIeHUiF9OxUkFcelyVv83scFeSREjyT0HIwi+eN+kqhlIxOaGeZB0PH
jR5fd1pGCZGqepRF7RG192DxTB93UBHPEylW8dh76uYJJWbZ/bwlEkrErjyiir6a
wHjMjZ85OyU6d7tAQV/2fZSEPWVS/zucJcOiqNYVV4fwCGCxuk4OmFRBTCXVHzJF
rnMbUI9hqsMQ3dDMmK8nEyvOgpRTQBvJ4HUSYQ6V2eGIcOrhDUYvDX2qmvNZkiHs
aG70Kl3iZuBXrKgmGawbzkQGeq667gJ6EUnstQ2eJedKDIqD6WV6Wa6rCfdzdw7Q
5QYG2xlaS8K2M//nEmQzxvltOc6J81Cw547YgK1lstC1zWme1v7AtDoVaaHaED+f
xqd8hJR1i5zXXG0EW1cwHFMKFa04io2A9RkS/9syNuZDszt3vG8eU1kgTyVnNil0
RkNObQ0XUtWL5L6pAhvazD3eDC04WaSaN+kgmiceUI5zJCJXLz8wPMuXyzRrOnBM
uxTKTRPB0piYvaXfBUl0NVN42QqZFatIImvgkam1KAWtX0jJ8u7DljClBs1TsHDu
mtSBQpnxI4Xrm8brqMn8k205mDMZBet/2AnFY47ARmHNrxz3dOsZNHPK66PgKr5P
giQp4S6R+t1HNgIWNeA8cF4ZX/PEgbadMeDIF38neaja+jPyUCbMkO2Moes0ZeeV
vGWO65GIIY+xMEn6ayZaT6YVGTxyUXrHRWtnSPxxu6L6YqRDy3M4uBpyb1d73Fpo
t//Hm+Pno/FNG7NhifuCgzTipQA1bWO2pm6AZs34tEqU/bV1yLV4KSD7FwOegcoM
9YnshIRYCmjW61Vl85HmRuc8KNvtXf7e/XBInx+/Brlrh2X2PRu4M/Fi2thrJbk3
dqAr0u0g7yprTeUPErAcgy38rRe/qFZDUW3V1gGvq5Dgq4syvbQsslafuNpWdpK5
2xSP5En0JTNNW6sbl4B8v+a+MtrqJyLxNIgGtf7NPYMnwRnnBi7E1P82Z+vs4Kpf
l5r9OiBIgxnUJD/rbbv5F5nW5vIH8JE1E3rsqbVkrApUjyKUjWUO7pXkQlHcHzEN
q3NpNcHw62JhrQTpZnq7wWZuNthqPORQ5miA9/2pY3iakO90cfbvk/psJU0XfPoU
wnHpwzQkPbL7k6MdrpgnqXoPZ/heoOOSDYy6HCDkhzdBbvO+kpJuAqYBR7o4w1N8
QIIO8OYN5W+mIvtKcqygl+q90DnlXaWLL7cIXtzg0j59AksA8a1Bn4qslu2FpyVO
jXgYZt8J6nqK6iIW5Yo6RGPz+dPkwin5RJV0VEzN1QEG1k3TJ1nX4Yrgt/tTuqhF
uoUTBMkz4t/aSjqEpnhdrL/p9Cq82OWDw8MRfSD5mJllSAE4Zg3Avy0L6h0o+roy
WSWrEAdb2qHUccx+3ZUS05RuV2iwKDbBi7nieONeS1f0L5BuoShUK7vAfG359yTb
gnbtzOgM1IacKAAxo9DRDKbMOPkQS6pBC1EO1U7FJa+Disg0dK0Wtvj+jVCceQwn
P5qbl6m4rursRKkjSY3kxV3IWzhqNLx0+0EmxN90+Swg0qqkXBEPoIWRuvTfGfDF
L1uC99ePqLtJM58Lx0Ltg5wcRtUtSSr7xGhAjxJyaviHBu/+jS2s6D/8o+cnV9o5
k8kREz+mX6mGbolK5JfL9FKwLJ6u+fOWYPKC1Ie4YZcy5vJdmNIQvOo1lXhi204Y
aBNS3gp0cXldKXS50w8BcTk435hoffbITPeAcRhh/clgmeeTwaIZsiXnMOnzXrD9
SwMMMOMxScPHj6dhyiqmD2Xq9j1n4uujoF2C+9KLg6vy/urmPT5kBEULXTRZWljg
gkomG1IMugBeQ1+vd6GfTvYvkQt9tvlI1fBaQCJbqxpA0tCdSZs5eMsf66i1w8WT
K6DkDv6cswY7zyzYCb1FYZidbZjEnVByiyMC/3WDd64iu9W2fU2w0TSpybLJFEdt
zrLOl7t/SQwhvPdzaTuBhdEIye+f8QwWwFuvHe1MgYFXSoeTPESNEvfnhi2rJGqu
BVlKIHYd7tFXfM5zGPmLXWF0BpQl/52kuDFLSHLA/+AD38weli/HbWUVa47eEZ+L
frEUFzuXVC339oKwv5X5Jsv+vAaBVHI5oGdIu7Yo2JmBkZZeHVe/GHQuiv9FO2+D
2GwDbMlqG3RidaA6JBwIpf9rU3UkAE+9bmIkZ9DlMGZ4wlyODs7+QRtC51f1ws+/
AI/wSH+KAEShVCV9Cv6V59PT25mxoUy7HkZ1uoO+OdCQZLFFI+afIKFvzlYxrNDR
gum9yKfPQ08imyENsxwvM98a5pGl67xElUYgJaFO+dnJk0W5c3vm/jimj+V0z54F
+G7G8h55j+eTZpQnHK3tRm8W2Zp6zqnx2hbKntnHchhDJ+VeqrU0MJ+PHVZebAuc
jip2F59CqwJ7wLIsYuHcNun5MhMATnD07F5QNJPJ87Jci5hojpFqbqYVLsEQFFws
vpe0nFpDZB1t/Tq/a//rJ5iMPjMuzhhj88dS++w/4Ow54e9zfwArjSssrsxWxxev
xEz8x1mR0nLCQPuD0CNcYH9FQHtQkLVVyIBtcM4xs+Mjv9rVMI2iBwYPLzEcWgxQ
XASFVrp1vQ9Pwp5yqhSXjf7HDcb6TFLSat8IFoIuER6yQr6Zr9b37BF9r42D4aHX
cr6zDk3Rk9hTtZ3ALH3hoX3JeRsH1pvK2ns49QRAP2V+5DcIBQ7xdGbQKQz4VhkA
/EF3yNxdU0kY4nYoa7hPC4NvdtTtSStvSfz9e/XtT+84ZKcmhGuXC0+9TeEGZRJK
WcRFREy9fhE+x7F2C6R1Md8rGFs7rGmvMS2BJSWNZOSF6O0bYO88do+WoegSBD1a
yT1DpYuJDq+c0ZBT06QVq1Q5wS/48qoW6KouLHx07HtG0Z+1KJotlY2PhrHa0UMI
JcDAZ22KSkYvBHYdiABXcR9LYSboxpe2Ei3MkUfcIXxxT07giRnWlpIvDJA3rz1X
bZFmzsCxTGolRap6ZQmwhhkB7Ak5KWS0TM6H1o0BCnP1y4XiwIFTauOY+3Tzu25D
F5Se8d2RHDsPUwMJZA7MN8CgGt53EAezdmZO9SQgZxObYjVbAZ7jXFE8+15c3CmJ
uGnN3qlncAUpYQ0MJiAnpQXfvwH+C23t9oQf7NKX4emhIUxa5CLucsHyzk/hmJO3
N3rGzGVm6IPjszSazRIy5XHHx+O/SHXEtXY9BuWfkhHQKkCDS0tEdnUhxeHsiWW0
5sUVBmlygkVhGqL7nQkpz8pTB7y0qNNd4Wc/m9Nfjcf2LHaVtBdH1WHZK1TiFroy
sZhBPi3JkShhMYTixgME4UmCNW7gkdZAV8UMZcRyQM7tvOvwCczldRfZPQAjdjTo
KI4x1WaJkLL1O2t0U2YVnQOPv77aHq9Vg30idbF9p4imzI8XK+3otJf6dzuUSO6G
kzO0fW5iU6aJYgmXYGk8Q5aAvur+I0zYcSZK+3Y1x6tB04mD1dWoN015mR96KYu7
ObMXc5owP9jm16HVCKAAtMZkvFUi4KPRPoIp2xQ3t8efNSnXFQA/cZPxVEunDFrg
m47/gO4GT07b6PoMlpGxzW/7WQw0L7VDd2LeZZ4qiaHKHxbJAitO9C09r7g/LY4n
aCA3qy8t3C5w5+EuKNWVKvJqavbJZefchd6jFVyoU+aj+pLjWOzi8Ndd3nJB/BOV
xyHxnHeWYpACy0O3RIlNb7ddOk4FN4i1/6xu+dnHoHvLeqcoyH8KF/qiZCsU5YYL
+HhJ/lPgEE3dbhnowVjtVUbib2kpGAnNj8gyYuFrV5h0g80SSxLKDUA1U1G0qnFg
dwwV5g8oM1D/N9gyCKFnsdm3sxNlwctJsa3zK76KLJ1Ai8v9Odgk2/7Sj55jrZmh
+duX2uv+qG+rq3iJwVBjHv1vz6jlJTdVqQAMWF3X8XFgg2nQm3d/vJpIQpipyY5I
bEWVCNiNXYIgXcFG3luYh7EtVp4qBdpRkOsReENYZs/8jSxvA/yS/vNo5roEDPjQ
D+tlskNi1MJxjJuEh4XslAw7KIGClrUc+NOkFCkEPjKapRtd5DC9y8RQ3fuWMWdJ
KXwabrXlkdju2rLvDlys+AvjUuCptVwR04fLdb162pQb1DjLKQLjwy1GRbU7XUGZ
BoRbJQGYuAtFdFMJpvqTestyaCcu7bl9O1lXoOVivx+YSJrwprAGpXlsICmbqR/2
ShYpNFn6GtQKP8LCX3E54KIN516VsgWfcdQWyPZwYqRqPjcKEkDcejF3HIXQqZR1
vQqu1clZJxK8ekTRhKWKamjX90DMyP+21QenwVT44Kw55JLamZzmmBZgc7YNKsXc
nKt56oTzi+3UR+yXlZa+Rxqc5VQuA+rvBxWdTgCTtple6jQbLv6H50giYFCCLGGL
ZYh8467gWa6IZx0FpPLtccLdxSC2JBA6BBC8QLl4idaJDmE0PYqN8sneJW8zUFes
Zn8Zcdr3nOVtSrZs5oz0a9B9tDcXDCsYPnBs5+8zpq1Ti8vscGNDbouaVhsYFSGZ
6B4LEjUfYAPN9CJPJ9ed31lPwF8sz3owBh/1AsSh0GbuGXUKm4PTWeIyc1UwMVB+
t1S6DcwUdQsYf2HzcnOmM4B4AiQyAYKHdimDmy2GLrA/fnLz1P2+4Y5ZgQMDlSd6
1NfTe6pQqndk1B5zPdsXYebyneb1FWJZPAlxniz50dcOt2nG9IPkzoR0lbcNys/7
gajr7s4dMF3yf4pFF2CqOaw/eNe9+Rb8U3cfLykiBxgWflvjLBQ+r56QZ2MsIXiC
B9P7vkQdvICR65mKc3MwpiivBVVbhz3+4bF28Z2+l+gQwWkbWAvDViHu8yw/37pw
7yJqQAiltdNlQewGQgsUIdiB5Tjj9rYpfGYEVntydUTbFxnyE16tG0qc2UCIb3Gc
asNGP12dKUZjXD4t8HPxUw9mOV1nXMlXrilstnbsnoqbZW74AyCLikmNZxb7MfpC
iCHFA1ZYrJ71Olco9JpPoOWUwCeD74Hh4qjElkhB27h6NzQjTu0Ea3/u3XfxknMN
/afIL1ehyaVloOL7e2LOnhEc3X/BzSoaNceaGCs/dHuql2Z7QXrG0gNI21kU6Wqz
m8l/iylC/wNO8umROCCp53cSVQ6pCHkjVBUQiCQOEYoOyb7fFY2fFSKza8SDKt1r
htGPLuPHjqvL9cj63qAsUakNCSfLm87rVT42vrfv+049vrajhppfdw+lQ4QPfX7y
l4sN/vRng3G0sxlqYC3fyVwHx1l8x2OE6Ks+V5A46oF7s5265g4ZDoycNk+nmjxs
6G5HdxahK5rsStmZswWZcWp+2JSFXlG5tbdJRnFkVepjVv3G5rEXs74JSxTN6o4l
oc+SNr/tJwN9QnoBEERvZMCo4aQMvYBCYLfZLXmj0XmlXZ1ZBTjjnoyKM/ubP3uV
m2lBPg30jMrhMkQh/TaIVKoOefeT8hyKt/NypqgPR2VOqasEZ4pi3yJCcpBGivr2
liOgox19mx+v/dJpzC2Dipj5IWgl31B1PvPljLETwXPpCeoEo5Ih+cVkcmEw6J+N
/TQfjRat4O4K0ysGSouEt2WmSzK8Pgicu/Op4B5Y37CeOBWZ3gls9hvgavTq/Fh8
iOt7dkrzbLal8l3rUUA1MAI+/4dMdnxZxqqmL0RQkUQ+sMNyurArYzQS1lA4/7JG
bOG4q3VgEDDaOGncratnO668F5RjbKxxua3g018bROtWwjF19AitHfdgOTxfvRol
z3v68jpYWrwi6Cr7vJWtg0pIZWJoUj2rvWiRLqWjLB84ImnzcuVSy1RICJzG3NFh
/AaPicNU7JkyEV77X8JPlk4gwBZUoxyaYF/mr/X0qquuFBZMKZftPcwNn+T53pZm
Z7S8NxyVfnvjmSUm2BfA9NFGbMSbhN7J4A3FKsxQCH4iDsKycYKoy3ZnQGeLqDEC
XGaqrHG7SOeoxNnptL6R+3XuzaIvzCWnidVIp4y4Tr35tIKQhJ5aN+A4N4EyYNsV
XzOWaDqSliW1KfSGLosYvkD0F4FiZ36ZyGrsbnZ6f06QJeJt2yJlwABb7zuCL/mD
qLal3o1KHeQ7TjdzYfMoM3WcBPVY56EKmEijHsnlqM7KIw/haI4EQBsjied79A4o
RkHvuLGZvPS6kD0iEk3Q0cb7wBO+XhY4Z1N4qeeQSySsF64oKw8IZgF6DqoRLWEm
W/eTgEEHbKz6M9kNNjwZLOWmxbYjYLR3uP1dFKC4gTizZ1Ywc5rfQZ+9wdy1TCiX
yWHq9ey/rCoFCc2VelcVLf8tcHa5UzOrDpKFheYJAGu4aJUEOgFNeVaTglptjJOR
xnm9syaR6Yw1HqJnufT4c7McwEQqxuvQ7GziyzVhqDENUy7H0DeFkxI92Z7mXZK+
42ZXpSeF1cfG3QlsY9Wy5HUZI2X5gHzktF9pgWpumutfjleRwLJa4qxi31hJrntE
h51SUjZE55Yl81RsWY2vcHIVzpVP9bVRxFaqb5+jD5prwsAAAv5YM1Bmam0OpVTD
YHLplqL9G93zSQQxgCR+tDv29i6nfzH1GEVeecjLeXqi4cWbMXx29RwiwoURMeJa
IbMZQ0ZGOyL7F77V+LKh2TLajnRtNFP/pfZU3PEwc49DlY733sMj6pUoO5y72ycM
NZj7ocqplRZ4WzYcgxrJ0PlMoFZSgjgGWcixtq3UBsZ8glVCITBGUwhc3DiTuID0
C9jgMuK+OCbzBNZtFL0zWnvj4c6O7eMLQnrFCzymbRxHtddDga1uXPIRitN5ltmR
GtYKHlKRYGXpAHjjGsNRjdda0Qmas/5reaunJBmj9czeujGeCRHgZ5UcYYS9GKFD
m7PrK03MpUn/Z6iVBWUo22ALwTQTlgYO7OsgTT0TqIjyOCOB6ZAMynv43bL6WnY4
MqQuvmDzSCgxhGIVIYssOmSSmHjx/k2cJ/osijMOplWOfQZ8ny+DTcRPoWSfSMEy
7qJ/O/cKYlebXVCW2kqQBBd/mAlF3w315sgr04NR4nn7ivMdMl9O2lmRYDTWtNtQ
XYRSRX3wiB5URZz25fGLrZVcuVNllQQ+2rQL9gvSAQU0OWV4ezEGa9fNaq4T58f9
4a9AA9th8knt0Zl9Ds38cTIfHTJ07L67byk++BPBmaLVH/6boLw3lMmxNYRw4KOG
pt0VWYB0lUy5HAPuen/aBzWHoBsgGWoiwAEhfPCPpwbscyqjY3BLsDjRmH1oQNBS
q0y998PsOo/dI22m8h9iswfWja5V9zXjamy9fHf1V5de18EJJeZu00G4TC/LQ4wU
CkwkIhxNBdtdbSpGOrG7AE22izUfafHt8fB4okZcAm2RSEcWo/8SbCTvJQ+5FztF
vCvxwjKKwAfVudeUFSOBhss+JeXv2XeES1K71B8jBvomKh715pQmtMPF0Gzw2h71
YTEWGXxNoTAQSEAbbVcH1pMsCWauewOrvaX4y9FM4cU+4RIp3LEyo9L1ish+GRJ7
LLWmAxqO2vBtB9tJbIxpe/XYuRuEGwU5KwG8A0+FxAHH7irwOXzdWOqyQULENDRl
LsBxBmad7ZEKLLIckxfAlLQC4uheeYzJp+5GmNqBfazjhWtqTw6aq//vkl37oDLl
EEGC+DESuJFiHhHeou3aJpQFK6ayRLAmGcAyNfJjPt1gpKHJkd50QZs26V7EDh8y
abTWq9uCXjG0Ldu4oh+xgt4szjVNfDXbQPFjreTkspikjYKF+/tfWQqzy7y1GakC
4lC7G2puDjFZBuyXuTPAJFdD2gXQCzMB2sglxpOPhsT8Wq4tumwV+wWRxsHqj4J+
QhyaHV3ok6ZQUvV3RNAbyx3llUGITbIv7YFI9ncthva6eFngF0ATDL4XSAPCJZzO
S1sYIfKtAtMbmEbcULBLD1EhcpdMShGK4YjgaORtvXLaCyIUNFzZRapkqFEXBZXp
GdLgsU1F9zuLVA+EK8Hbbufbpuw5VtngEVui60Y9YJNCgkUiZJGX8rbrIaKws7g4
hhN1oJ9Tiywin0DYRRvo0InzhQI0B19Ae++PSgXBY26LgFm9loGhTjtdCc3nD+XK
8wKAf1w71FBvtXnL2pU5eNhsk8AnYAZ9pWEghGWVAkXgb5f7R4rMXbMFNxvMfCa4
pHEROeKFdOYY7FvB8Aw6IUrnyBYySWuV09UqnfW2VgwI+MJVQp+IQ5gSJQc4S3gD
UEenbSUue2oPNwkIJiBzhenVAs6mpRffcqkWVFVR/WpclvFIbplY/cGBgp1YlL9a
v+d9WTqfPT//r90wQC8209KV9k5UY6kWDMWS2NvDZvYMu2TIvDgpu1qKN2qbiOfT
emrUf50NVSMW+IuCTMIVDqG7bN/ufsGzTBd0od0k4ENKBjos0qvO3kUvTsCGtgM8
adogDiarQbQrt8oZn9dfLiOAuTF+ARyLY7WZkqQ0CQpEm3+pq6AgrEIE70PcRzlR
wMsh9vmg44S6WZNryAt4mD1IAa0y1T0paEKVjigB9HXf8+yTaWOo5+upZSCBSCCC
vSJyIVKo5fkn9/CNLf1ZCySIeENmTDd1X6PgPeM3zIVGjzYkv0MJ5Yi5rPpLo3J0
jG+n4btSXDwLFcPm+eu3Tz9L146eyAHuht1bWFXmcCucthi6apjB2uZuzL4lIejI
QAJ63etgY0uD12Cxh6RVydbBmNAammeB4WqMtDhPV4t3vDJ8aqOoeVdR9wfRLYCT
zFXIeMH9+7N3wHvoI63J7jKn7bjstutW5El1izb5vBE1mrcq7lhN1c0coUule1qR
gsQt8p0IEsHjfk6I6jzNtSg+3RAbvI8s3agNgoVWXnYmSr8fas0AA4JJ/o6gyEuZ
uG072dvXAumPLmTVA7WEJCXrI0+whukbhmt5Sl2ArJIJ5FWkpd4p7ibPg9AaTfej
iTaN1IEOvg1j8GQTICD+WPpKHTJhKBcvANtkKvzgc8Gsom4X03SlPxr4D++qltpq
pCCzztYXDoSH8Vli3O18h4PncpseRptw+Oz4pnMAPC9yHK58lsCOTREPiAthAKKg
GeRYhSF5W54pyforOmrNPNB2rCP/PMC7e0biWDIOB+6DCBvxeEh72FwsZEwaERYf
C0EaUP1rSmvn0LycDBY9s9n5AY9TW8yuSQb1+t1cX43aW/O8asPao/uQ7PvSPPp6
zeUS094m6ijwHSqfAYCwvRnctcwsmllbebTyCTikrILBcwqQBx8UJiKmh/c8RaAf
qpOKIuq5+/+YHtOYcX6SOv/b/OY3kydKi5VqSoQ+BFB4B3a/ssZT4XRMQjb1vtD4
tSXavdlhIOjdF9PdBlzmCkWZkHbFqqCWjbS6Nb8TIpuXLXSD27VhpiqYMufF0qhi
x+r3ru/Ngy9FEi7wJPCJS3OkZwWC7fPTc0fwygQpM3Bb7ACFlN54eh2H0djYWNdz
vDasyrb2vx2PmMu3yd6b8CTmx/ItQHrB8ayosVvbGj3zUhDJbxifqxUB5auTiM0v
W6ODrqWSIepk9mzcbLTXvFe6tJsUnd8Fhimp3UdkXzvQrt6TuLhRaipWWzhpz9bD
I7I8XduFD1ulQBfn62X9iU2lHAa1SNPVak7266RXl0JwPQWg5cXzEdY+/DRMj8Bo
TSycBd6GP/MSaEhRfL/Nv428S7kOVVrjxSdd2fchMO+EamKiGKIG+fO1ZY95tplj
VwbRziM2wVeqDqxTYuNkhVBH9OSRjITVm9pr7xQjfZMbdMZNS19lieItbzMhTOr2
yHa5MJQ70JJl1hLl1OaukTam5ya4Y4Gtu5rjyfOqQjc/CmtfwPK/r7Grb7mIsm3W
ZCGixbIzgDFqKxe1T5KS28U+WSaanVpBeu0I87r6IHczpt1mQfXSTvoymsTu70pi
6u8G4VQsd5yTQxKmTn3ND2vGN7Yx/Z8HS4xfRu1XZN98rBhAnGb/zMlU1tCPP7A7
CaMXrCIg9VRaSdnEkYPvauZgkmj3aHW8I7qRhVo/51NhJFx2EhmbAe02Wf+S9HWt
tXvF2M3iu7nBXPlcECX1uv9HGvHUknQpWVKi9GqhGcdBlyMXo7z6VorcPPImYEiX
clthmqOYysfTDbo8eNB8Nvgi58QTVee4f5Z281puOASyn+/Y1VCTiRtBDSt4/M9G
+s2g58M5gunFNkjC3pz+MBBfW8wbRYN5zrmPC8OxXhW6vmhO8LGCH0EFbVRDeRF6
fV/QjiGcA/Z7xu/SSs+OleNKu7IS1gf76yb8zfQPBNv/8w5LdwMDOQqIN8nFUBMH
WnYdJL38UvYuIvRpAk35WdCyR6IgiKL6w6pVzswkEs04CjDUYYHZ6Q6L5hd37L/R
j0jp+zhf3TPxW72Y4dMqmRMfSoEO3Jaluj1aHETSvvyQ3cOfmGnzzI4j6qUhIh7d
efq/lHOLGTWhxmeBOooq9vT25yauH3dxGIOrla0TT335ttYBr8+NVlLDk2HkihOP
Kb4lLuYuFlRnqCQN9iPMde4u/nT2JLDeNTy/SXFdVeC676YiKdN/w3yBKC2Um+/s
PiYlWWUBOIp5qlQv6bS7CwGE+E7XG73Zb+5wjKHttykAjsJrMgFDqIHeUxRKNw5g
hg0oesS7Q+4Efsl2XB28tnYJYqwphYevaa/P9nm5DycxFK+oI67Fk7pbhvdeCeA/
F/xjqnHRTdA6nj4Z14OuG/M9tj4EaTHA6xqFIiN5PD5vgF8W+YeXAcAL/GDnNUEk
P3grPygjerbXZbRuUIswzzxLYmFEs1WLUI74X2OFWvevmV1WlpHtHoI2tUqowBO6
makf9nr9x8uYRpcoufvDeT44ObK8KNBuK8YPFEDTofSCmm3T54eJaFYsY1Z+cpC+
tigBGSlRcrqvrPfSEoT1B2zLnmB7iYJojujMGk1wOVMNjv21XSllQ3tb5qnzBza7
W+mbK8P5sSwcgB26jNETla6MwB6kWjrI3IiM7FXOxqbr02HWbjfiqmabLDsG8dIi
P0wJ+yqcaH2pqzI+WGoF+7rJrBWIkN4ta/l62LKfZAnHaDLt/w3eiuh9srn2CdtP
n0dawt9fk6xtHb5WRJBZc/dgCjPUaWFc82RSzctcHE4M5Zcp5m63ymVj8bgxv3Wx
+UFNObAjz7UJ8eZozD2iyB4QkOrHOdvbhxzDzq8tCAgbrW1MrHYcr7MA69TsrQxb
VGzA1tco2NqvCJ8GWTvXV2bm33eSm+EjPxOky+iprGquX/vicnj5xbPOQjf9SD+w
5eVqa8DgV8HNYKWXWVUm9uyL19jnJK/eSZJAq2WW62YKgpNkAfchTF0BjMFEDC3L
GjQhn5mlS6G6UNUb+8/342Nk1I9uB/T6iMvOGwvv7LtyO3ErHRaGWNA7fgRhme2l
8tujvvlgi5Rdu6WbdZkITkkUrwOTv6wqPkKAnRdtbhs57O8JBnKqzlHg8bgff7wF
aeVF+6rZl1ZVC+LYm7un0mTYx+rYs+tDU1raOw2DEWjLdKhvv56FphIfRxPfPKsS
1MLF2HbLrQjD2c9n0nFCvbRav62SPNZ9pABj4/RHdOWV/ELVTpq4SHDdier4OnEa
FEQmstN2RAEQ+11NDFd0oditm0etAP4R4yQwS2SEzMWOR0bdNKxxidWgfpbaaoHo
357y1gk/IYp8fw49nPkQxR3EcJKck7OuOoaluymk57YFoFTKjccmAsVG7dzSnBpC
VuaSTHjp0o9r+rzhggQ8Nhp8UkGw1//OAtelNdulsIsJrp23wTSyIlj5vbLZSSMK
X+Yg+5cyjExMUSMyExnwsMHR3Fu9ToHcKLsQeNdIC4XoaPnn0QrESdmomJ4rbV+t
hUCumSURFQ2DQhwuRIaoonKLATN8s4bKLPJwz6Q0fB9OCinfBOk0ydWEXvDCYxm1
Z4ir8Epy8Hhlpq+fyJmHNi7FILCVeBGQQeIP4Jye+rlGaitE+dZk2VHQSTyk74TC
axXBPTQx2g6i23Wpq9GXj/OfAb3NBZLR38/Cgk8IMwucKiq67OGOY0xo/iHyjno3
xe2SLW72vgddAAG7jI1vqwFT4hIt9W95EYT73vR2CP9PytRMKhBZXJNt/STVIGgh
aX9vwwRtK2PO49NilLEVSef8MWszjtBqa7UtFq7NPeDK1DAdF8C9TEIgBP2hZg9f
LcfjZmJ8/bHLL5+uCwjHSbtQVuqGMCOmjCZilXE7vnIKx9gmMLhaZVcr2f9dKvHN
ZAyPJo0Hozl76oxYSVrAJ2cX7RA6VZhu+G/C1RG7qITCxGKxNnN3EYW39kUF1ICH
xrzU3KJy4FUzQf8Fg/fr6U+JSWQIV298lmayfuzPKhvsItpTHu0ipFlWwvoK9qEj
/vFmN1v4My9ZaQTalBwGT2Tk6Lr0/tUPAQBP6GPHXuyBRnVROD2Puyt0fnMIbJIw
GMhOPVRJUiiL8wwLttptW9yA3TOlUzbm6vQtb805qp1/+go3ezv64uA4vDseWhit
mB2npqVik/carABDr47cCYBA62Lrz6tIz/kipbii3ETJYkXBuEX7x0FqaWjPMIwA
KLbF5CHEC1SJTR5oNEoh7enZxdp46aArDlsqX+mCf959kwoiXMftlVmgt4UGGo04
27ahbCNkd93bqOmQlovhZQXZ/XJS9JaAy+k5vL1HJ8/H7GNeqPyorcM6qH8dolfz
kJyGJIdKfClc45ZIMEb7zMReMT7dx+aCMbMPLoDG8jfqMqlSxF/9obb0syiBRfih
sECoT/Uybq1ak8PN/XJNBeEY1hT1TJIyXdt3vUUQI38vaoWsP9PzJ2eBKF8WLBES
K7JO3NFBCP05NemKc7wfsD7JGVReFfKQHOJpKrMnEYemDMPOD0BMjdXMiVY0J3Rw
jgAnDzXEgPc9hgRXkdreRZlyYuG1+mSjFWl/NMAFAxb+KuYZkrSz9Jv0nTu1psIn
0i5xUa/jaEyqZew88j96zwzXhwBZA1Dq0qVgSY4nbnl7FoGE0zFqHX5Q8QhUfdK5
6KIEUORF82SteXWVhuiEs7ZfvGlXKlGnj0SId5oJYIUubz20Gt+ThwhqowshWZGJ
Ij+jsPDC30oKLKObEAl9c61sKVptZF9sszEimboZizkDXRDn58d+XhpLlZ6HPB54
bKPsCiNBXkvc9/cP9v1h53z46X3qVNEXVM8m27nuGXV9KLY9GV4PUtMHxUD5GarV
xxCqpCZ1pvtyMljQ5ntm2KtbHvBKN7F0UE/QLhOnVeG9+maF588qzBWDUjfg2k5b
xp9slU3YEJFlQTayvBD8Ux91smgPHSF5nTgy3nQXGEJmpSeTrREj5w+F/TY7E74E
dpi3UCh6okfPAxzVItbpR4A8KilAixyfrsw3lZJNhiOj3nbAv7Ivv+ObYRTsH5nc
E3j82udrbV8vZ8KGByl/7hKVix39qiGqisyuuVhsN7rZ5zZWm9frseGMFVC5BDpZ
Fh+qvTyQ7VUWMnYr8yaSv+HDQ6KTQV2GyU9qK5wClMwGXIFtiOmMIK/adOsg2tEV
xwea+y2gAKh/E5Lvd8qm4N1/6GLNQzUdvzb1hup/ARzTvMsmZNYxj6F7QfzmrfUJ
YuNMcIPpHnAukSixtr4AzXu8Yn8LdLOb+IUqypSm96SnJoaxVrwdz6K7Or6ehXKh
6N+NSNuTwvhGaoQHPP8rskUjzw1N6iC9C/Jsyw3Ei9UhKrYDz6VzbRQAlSiXZy17
qNK2NvAlnHQynCuY4udp9mg6cfL5q9cdgymeYHdt1G9980C2TI4yls7t/tAVMRhS
N5On9Pgl/2RtUhOo5YYCURCuf8n983UwoAPDQwYAiuw7yWca9VsUiZxMHNVC8Mix
S6OaPSfuagehtO+wyWOblkofLSsuu0veYKPMqv+SoTulBRV/aCKpT40G5gOE1TFo
VQg4wWDsIvm7me59WByEHIapsff7K/yaV98nTsUf96m5WdHypP2eJlDxMGHyaVf/
JMZjMPK4l2p8cElGLJPjndD/tiRn6pBoYFNXg7VQ6OcuwNCIuUz3phsHQ0yO62SC
Dce6ZMUmawxQYdE8B5LR2qLK5odiQ2wSYoevqFzM0smECl1cQPH9BI50hPxnHzzB
kPX8mPbacSyN/KhfJBsCJQatcrj8yWzwrJJgoAsa+bmr9Q/QuXl6oqENsMBv5qeo
T3yYY9plUw22k6n5q89ql4kkWZVu6F53miN+RUHDKD63ISCTMS5Z0QE6arcY4dz+
Ml3DUnXUAFFLNsiFvrig5b0t23G/RzT+hg2freLbQA15D6Og325VvBJItzVXuoxc
Fpp4Pyq2vjls6MexOHUl2VJ2jrKCx8DqbuOyXCbKAwhR2ZeHwNQzuH8U1vuMMsTj
NPTSgqlWfhyjN4t7te9gTtlpS2gkoOh6J4wmExCSU3sHo7pxMfPgI8zNo5o+sOtj
lo7DULKmf/+OgRdzcqwz6lszOG64o6hn9eX6D45HuDTpWZjoTYrPQtWbVRvu/iub
j0mhbH5vIverykpqxFJqWYNBDNKM9Axh7PCQe0QP8JFEeNeV7A6ZZfHxYAdl096O
JiGKKdcGcDtzMHDIX87iJ6UKJi7NSGwQkcbRtHRmGlxSMJ8lCeZesI/3jm5I/Boz
dkXdsC6Rd8Ao9S8/oDMGLGF3GdI/PVbmBpHCjXHKhAh1xrYYtheFMILLpVNHOQ4m
l0Xbwk4krn8+uCtg+7gYgR2rEMgpqI9PwCbL1figZ9qaamsjuQUFskbu2vw+9CTT
SYz5kLhNn6XnDBrl5TzK1UajXyMpaMlv65nOHhrDVh/eIwiTrJRqGyumAmxI+yYj
xmRnHzjiZpo2oCc8aW5mFV5rwicPEI+omBlV65Xg5zJ0WRUvELbQUyOcZq1+YdIM
KP3stNWmapZKhYGt8olBlLsFHNwNs1DibfmPGXEFLevsC8ZR7UAC/ZAEtNroairX
xvoV6HCUpYpZ1dJ7SYv7jp+1liXkiFFyvEv+0R0/3lEkjY4IRPLEEchKmGdTRE7J
TO4rDUYquFEU7wTK4xg2rNMyfj+wYoj0Osy440xqWRnUoINKUumKgS6Eo/TkHzTA
0vYDmCa76bzB0XtG7EPudGbm2gS3NNZESRUbeC/l6AX/3qJkD1Vhl9i89BG5VJuu
nfC1kK+z6wkrpuCO9JwfTz7d3RDK3OuwOVa/MvLytxISvoZLbkyVBMBM8XBX3W45
Z4/r6BQjVWwSqLcuYkWueIgE5cvexCZCQ7lyI/6WsyVuUi+kujReOnMxsabUaJy5
xnM26dj1sEkrTP/8zVUvyRgDEQ/m/5WLqDHB3vMfHnZyE/azEQYUyM8s/eujR4pB
4tNB+fVpF2Ts2LwoJWEfHfxwr6PD1z1+npNeq6l/Qkoe3suCRw3uOQgn89+SnFO6
QSoCqwMoZxMQ7fSJvqykIlVfsduFyv+9D5LaT2O4D96sHMFt6DLCEX/m8pDA3cOI
ICbo+nz1xZkXAUx/qX7RIiKbjq9kFBL/zQDIX/YmNLKNhrftplptwouwKuZB/B6Z
Pfw9zyMj9YJXKzwXxBJbZtmI78OZuSz7jdyE8S1WcY/gxkYdvwK7gYyWM50wY7ui
CmQUx3U4yTGCkZIuNNMwYtwhQwuPTCrCu4R0WVa6FqAsKPASVM4+2FaVXeYXsOYU
gHvnZCCWuJP//gTcBJgmk1juMTnOlkJ/k2rh4Nclk5Mra1LhoW87nzVDo7NOTfIS
k0uzW9M/XrFMMD44YXSPql1I3GCKX1E8elnhKgk7Ix9CQWSIqkK8+VLtLmn/uy1a
088bJ2xQNdjEoGS7LSr9IkkE3XQpdwyuk5Mbw3QPDf/sR4FtscDWNZ0J/CJvyZxn
bvluOIm6Znx/kQzAIdeHRW6YhK0p/Mc3atPrVExxBcMJK+mNcvzXgfqUBK6rxvQ6
TyC2ZFhL8xRfpDliv3YGWJSXi18t6gFPnSe49e/io0gNLJghhsPr9ttUujdsDFE0
h6FrOMIAuntv4JzwWd9dYQujeewy6g+dG2a2CtLohEDP3FY9Z+WtBMorNfhCFhE1
PlTqA1c7Q98b4CTZu3oxYpzCUDI7OXqVtD0T6rUV5c1ac6v93iTNEyIZXrYV0LXZ
SO+7psXOCvRBqKjQ90UfTmxHbtqu3+r5cDUPxb13Y4JXCRy2+H9FUSTIH3poduAA
1CTG/hT3b/NxOndfolPDVt4smsY9NhO0KW9z9f8b0ZCoUcotPcwmeXM+GSy+J1ju
lLmnFZiC+0zu5fCJw4AB1szc25uXpElGi9nm4mZ0ZrpQqsJgw+XU+AMdTZ6k4hKg
DRttHVhFLMusqsWYx1fd+11ETTvEHZ5TmGWzjM+OrU5da9oyfuauNOWozNbYYsNY
eyMZJJfPCmCCz6GPa8+BF/6GEKXA2rTwPFsiTinxz8p0vXvmvKKAsxO/RhVnbyys
O7o+sygeBQjRY8DYaDun9SEtQGzjS/1wZ6CkmBEWSfJmNrlNvJW2ERsW4TwWFVLr
uXSX+fkJjLzxYhEYovat9Lc5pY8m3jMMqvWEqhT7eUqoQQDotXg9qYIfy8P4sDHq
AX527c9iUgd60PENLWYXmSUYtrxJWqwKUmWyCqH7VkMIL7QhA6dFPzrAdKgWDI90
SGWW5lnm2gdz/wPtZp6WloMx5WMXwXPBxJgIkQMbsBfaYPD+AyCAhUCFJ/EkMQog
HWqCxRlSwF2vsDDuDNizLOBjlT7Wb4UIFYeD7glRDNfWltK+BdYQCeGjl8FY4lou
hp+CHvrI0KwWw76kSAjj9Tn5vGT0fVJZlBCmxZ5MbZdewZ6zhwCBRiIGh15puoXs
3cTnu48+oY3xV1uWlBnx/+sP7ry8+cd1flirMIpApv/zS2V2/OGGhxkLGr+H66RW
8qIBa0YYGDIvEmeOaes8uife8KcODVmc3jU0guGJRI9SPq5hP/3ZjbawRXhUxoXk
bqJ4KzhET5lqLrg8M+g4vckFj6M7zmkUTtKCEEMtWSmjYJfLg1GeOwQRhXoeXGsl
z95yt/0C4u7nAvxhY5jNB0uaHvgscnpaCMOR8Y1raCMVgpooQVahO+x5PDQ1tkuQ
Ba/D3rVXJTLEERZse3TwE4aV7BqZOvbVE7WDMAtdFGkJGRhzC6Yqg0XnKuw3rr/q
dwiABLyC0n1cxPKt3ArgQAppuI7JGTsYVXeII268Lyrq4iTKviwMsF/RNd57/Sov
FVWHNfI+pMPersQXtoDHn4/FlZ7+EAAM7ghTeKW74UFQppkGNcJreaIhdg09/Sep
rexfI2LBmMOECTjfYg/zmOR39le8nZJW8yNh0nSysz+Maqiu5puP9uUqbUxIOrNA
6+MhYb/mU+V3HsXktceEXqOGrWDlqvQk4KLULZQRc//CnNrFGWywWPhaHt8dOYTX
NCO2ACSMwC6pxKQQpspafLmVc44O3zsP6ZOITD2rjXWN+XE+8vw+fN5iB2tBAh9V
UIt6nGj3OydCp7y2Y8z81I/H8mBDOiBhH1tuKgiIeMvdHOWa/EsDUclnevkoYXte
CtL+uzY6O3SYRYWUJn5HaLlmwD/a+4LsHsAh9/gyF/bhdnYl5wc5EPolseato9rU
3B0tqM/6ipwhDzNAD0B62WL/dLNc5dIMu+xb4+ZU9RbflIUutl2a95345hnE/ika
mo/KfQXkfWmTMt5KaSsxei/VGJW4sGxuZSdOQN2NRftDCVYc/sqWSHd1H+ai81nn
XLcwGTRmZI/7JDdSOSJQ4W1DlOhhRwYNfCkACCw9nHXqXtUusunV0HWStdd5itG4
8+ddqFTGEDabC6XuCVOoIkxxr/i6QmZRhBqqc5+9oVa1gPfgVMCjaJn2nkpyvMN2
oqV+UHVCuFCmQcrN2wXmM5+hEZ2VGnfFTdqL4lBQ6XHKN9M6/kMnFlbkmP68nEPy
EKM7l95VAhhkdqkiPFyKhmPqBNI00FkfN3FGgYC3cAXmBzNGtM15rIjz8ZHW9oiU
SXW8No7u9vwgUe2U3GrfLonUMFmuimSRcPFbPIqvuVHyxZedTYOyeO+MRYtHMDgK
tXu/8/PFxFI3aEcvDTGr1ifyozFTfpYC1xMRhgiJtvaAc3iqK8SJT/msr5GPCH+7
1Wa4kmAYkpBwx4Su/tLIX2o6xq/96DilU0ye07STFvA/PxEXk1ib9m02m+/CXwMF
xSQKKDNZt+n0Tu/eRsLze4UMdNrgqv6H6zBgBkTIik1vTUQxEOQ4WNbxmMxD4cds
F/1R0AJijIhK48WoCv/t4Yz1LZYfcchT7QgqXscW0RGBVtyz5UDFpSl1tnB+5/gt
/jG67EyQnndxWZx2XLdDzxZM8h6TGmi/aP7eVjb6Ho2wofLUJqRCenYMfXqw3c0y
899BAiYWTG5psgy54zaDX2TBT7XhaHHnlQDlal23Fai0NzwiP/aLwq48sdhGETEg
DRPVEUoKn9rsGj8mqU/L+fJGrumFImXb3aRJ8tOH4RkokFMbbVYwAcV/TDCkaQi1
34SnGa8/ZqDBa8ZM2Z4273OetU6XQP7syKOqwy/jqNsGs8C7Ymof2ChTKjS5DTEM
OKGZ1OA+nDJZl6mGl7gOaWHjmkGkSwKBv0cZH1ZDxDuZ3uMs2l7Squ+y36qh5+SS
lhAFUbnglz9300a89kJrYKtV363ErWpjQ7aBTBr/jS7LCl9RpyzkYY56Rzx1SMqG
o/WHKOxM7jtHQSxDP+wuB1MI5VAbaPos8mzBYM+VbE07GaGKcyDv/7HDethpDwdy
+teavjAi7aQ0cXL8Ridt00BJCZT9xIoETa829e7XWeqQePqrEfsC5BevVXninsBR
aMm7A6Q7sWhqEkLi7YmSb8eUVvDXPm3b4BnfPn1aDmSFgWdCd4aYZfe75KvSyzRp
7GlPTHdPmEsKvrNT9Mn06nnck9JlUnrgIRRWAMA7KmuAm5w/tpgqMHw58uac1xME
8sJT4v5W8uxg4RMOsIAUu2J4ACKIu1CTbRVOlhl0y9gerC5YifPWB1aeN9W7IeZm
IyonlQG4snbliN5fK0OSxuAQhcLhnR9436EwUY1Yf66x7vdJjaBOHj1wbfEbtWpM
SlWUQyoIph4dpDJGTB0SR4N5f8gv+9axuk2JDtj6pFNKd8w4Ogs1U+gr6PxEoKqd
zK2XChydAzwD9fx6R+l8zv9iN8KnNkZcivnDAEecD5IbHQ8aCuEbd6uYnZ8BJvUk
5PnGPMmbVTb5LPeYI06eLxGAXUHIUPCCeIbJJbyKD+oszGp1ae2z5GSJjIqfEwM9
e0KDHZnDZTkfs8Nai2aQTE43L0+NY8epdKPmgUzKuq5CPbRngpuEgziG1uEr6Ixd
zXlELI0vOpAUCTyBdCQwUfroyoTfjIL/IL9AeZbzNveRBR6YTTn4vmAK9dYl+W2O
lChGO4e60/UCz213Qd58MGhP8A0kHzjH31SAWX0lkmXM/GPfvJQXSQ+4To0D724W
hxcntPaWZVysVInFl+qjxnvk0WR9lnFiFpegMkeoeqtR8BJxXIm6U6h2n0n/ve8G
1mvPkGEeL2hm79EnrDmWltEEWSPFyLPtc2EOf6eGufJIkN23MnRLIO4sVDmDfCxM
/F/keEaQQfdp3f01T9sof05tV9QBQ+670ET1bD9B05Qsx5jzCRX1m04WzKjeu7tC
3q7MizgYPeEmvD0722bLl7sxWQdpK4GUt1R6DamSh7AzSNzja/GaBIIeN0O3KobG
B8zJVmpjrYfFpPPH8WjL4g7GZTVeO4F2TexCdrtsV+3gs1HZLCkziqdetmtrv62c
C86qkWJAPGpQfNrlcDYupdWnjGD1eo1MYNKLhWiph4ZSRSehTVonHzKV+QmBGU0G
hGYGKeOLx0sO3a5LANfwhZvCrKP0+xepJKJNPKkXibvGFoAEElOi7lZLWJ3iM3C1
BCmJiWL7ljbVHdYfDVzHu2GyV9415GJYWkhuiaXnWbPdXF1yLkCrYlIBnmaOaUOC
s758VoXYCshc8FB0mkrdCb/V7LYtRGCiXwVaqyx7I84ajKqPTJHcCn1fJW1Sr8ao
/Z96tTZx6LyGiQDHULypXuEs5q5ffv8zSrkVW65QJjIrdYDVtSywi4vgHdWO6MhX
sVTA9PYu9jQ1AFYmYIb88clNm83b6dDWqlcCuSYraSIya3HxZtsq3DdY1tA5Xsrd
HsR6SqGtEjviLbbJ4s0P6SQ56brya2dlkwNwOZe3XpLsogkdE7QqXWmrUMeHBzvX
lq3V2dkOyubFh9VXSvAiS0iiFAvn4Sz8P7jsORh2R66Cg8yJbKJAJR7rUFzEZRYf
F9zr69L/60wZkGw449ottW17XUh49MHMjympbq39oTo7T1nY0P8E18KzdRCQIRNV
3ZyD2gspP91OtLiH1EtC0hV3QZ2IErOTcIpQdOFnB0nc/sZGslj6uKCQK/ZR8ILk
nIzxmztKTtHe+x14ulUg7URk3EdY8uH92WJknXo/uHQZtuhkh0O3xD8g7QqLx68Z
yLkgJw8PAiUnGQscZh2gzQcdgGXfLklICgPje6g++GIzd2mJI1sNluT+gM67muh5
OKXw4/56hy73EZBa5ZjlqA3aDKTqhSS1D79xvkQax0KjO1iNeaKtGTQ+oR/5tmKp
FamyWTd8KKYH/hDcYFq3yxmHP8CA25s3IHw0RM2DpU+xQTDWbQ1tBIrbB9u605h8
cgpYC8AHGT9FDu6NFqYWZU1sPKQiE/aM6UFlPYP9ortGMEnC1Yg05B4FpKEkAHP7
M4CvT83flBf91jg6zvaNY5CH8l1qH77/3SeNv7dtOoZb+v4WQ7TS+2AtvvvJbUWw
T0hA0mODgcajEgAhVnOxDMHj5VhMd8wlxI8qXHrT8csilxGnEO+0h7tIj+9PvgVh
kP05iYykufjjoa+dEN694ZMD6kXfmZIZbV6kukELB13IDD6AK/+0nPpTS3GtA/bf
+BWsPPhxcV8eNNDaVJtZKKuD4MR2+53bk2cEcelMxhGZiRl2qVwdPyJIcXpx5LnP
e6/ypIGQBJlaOMUx65JLFegAoUfUDflyf/vuCLhAmlGnfxcScCFVYJfuItn3IDUf
3n+3JUmBpI4QuiadpXe2ieiLwjsXy9IXyWs5IwGT+dGYrk+8/gn4A///6cEvKocc
B66ce7WcicjYvMmhYO0jc8kX8Eq/vpyrHXw+dN6jlNMZkHki44OJ1bHbSdBb45Ln
c/77Sg4KJZa4aTT3+Ze6x9zfWV6q+bYIM4W3ZOIijCHunE8VoGYCjllqipja1iIW
s6+ENfuswN3biWBnKNMv1gcTe5XV9PrFStozcwYngXHKLncUiJFAnpRQs1MUpkzj
w7DxzzALsC9p5+uVIAVTZZ1DwOrJj6Eju6YGraZmkulam510sJuBhjMzlmNb1lLl
gA2N5C5/DPVc7WhC94NARFlEY12XLd1EEFLnLWUNTks+q1DwnitZt0JPAo7IxagD
0FVXkldSXrhTXSH3Hc/6ZyQokiBgn9F1dCHwI3/QY7JxF4f7ahJ6IliztC9ibDmw
/vT+YoEHlw3M4+dvg47hEZdCPT1AkESuc38lE0K3sHZtS2hDguXfSNKFB9XuJvSG
GMa8GOhfpP3uw4DefHC85dMR8bEamZvHo7XJ2euL+sIMG2nXRP2ethZW5DbMO5q+
kTQCAYWPgM+OuCmCY4bL1moPp917B0HGN8RQ4cQOE0stdYRnPQUjsXH/acKog7OT
BW+AKZDtcpNRn1eosdQi6qLpCeECi1zzDDTg0Ix+vL2wlyaNsLgKDdGBSHw++X2P
wuf37EpDlM/eO/F38I3poswuRmDMXGWbvkiaUJLBfRinq/BnP86OKNWMW9j+mgHy
HRUZo7bz94MH/Y0+IthSJjpEIshp2bsvOgPTZ+TTEzoYQWyZAp1WI4kGuOAVnfmv
zSjf/w/aiWzHtVglp1NlfUmBvNC+tKSIYau1XO21cA1WTJ5rSvbmq99E2WZB3Alb
rFivqhE/aqQLUyt8ORHi/ivXhrE8DkB9331ssAF2qRDXM7lVMsrZuGBWM7M5s4Pw
/lhkdJ5dT/jTyKe/l+j8SlI10fjy0Mh75FHK2SnPYgTjDdDa/G1j09Qa8MYNX+jr
39uRUnc4gus6YWry0NUwlWtlKUwjJSv/3uzA8aZMT/zAucRZ9PZEBbP6xx+mqkZv
swJM1Mvre2ZbNAF4ePE/Q/RCrlbvan3T3Q7qdQj0Mxo3p6MfzsDEUnnNQ/oB9qAv
+Quqwamzke72uws8uGvbyTIFzvEbKL7JAuYQNugeBG8ce2XngYz/XUPj9XxboXXn
dBVIDvNwbROZmVat78MM5v+8cjsA9zNGjz1lpF/PDBK3+HFCwL5LGWNQeeUBCzcm
wDnERMbnVbLychraC25/g5SShlKARWC54bxxiNmbmMYReJOD5vCbMviaNHePqqAU
qZbC8UY5LhmPadJ0SEaMQ7jQcft7Ui2Rl2bTH/vRDaUVALnJVXhJ1TZBTZlTOjMt
CkeYe79QV6WGiie7c91fjyeloM4MoexQr60qobSGSo8do8pHjJtheX9kxMA5rbTd
f1O5kvrHeoffvv2AxYMvLx8BlhaaEaE/EJ1EUqeOaa7FkNXQ91iILaJU0/pkE3Mi
uooye42NnxyceTdwWwEShhf45LP0Jr28tQ7mGXrtAxSDrXqMInIWpDOud+6onTbV
41FYWRyf89gv7YOvbNBkKBJW/mOQk4rQBKIlk2/fDdG8HN8s/AjRC5P9U+UBgtKS
um+USE5+wGAI39IKCGHyEQePmHa6sxJLp05YPcV620sfOFneJjy7mM5qXnvCDPHX
cqlalktCAfTOZqSFb8l5cNNhdvinHFmZ/S4xLt5W7G8WXwKU1W//N8WbA1/F8xqx
11HYbs/9e7qO7nwEIvZoph5frU2BEGURY7Qq/dGL8avZTxlFIjrV2sIuunk5/5Z3
TW1964XbOPW0o0YIUjIdqRh8DPHiMq2b9K7NdzurW/zmblMuSDY1jn9bEaTFe14v
I1mNHJkC2NFrWgE+4LqTu4QjlCywTNhReWiwARtBBJYuaXBTjPe1YMw1BmmcCLUl
4GE3xAG1vBhXusiNQva1HRJJQQjnGvkUPee/W92NZHXLOqPmmZaH9tfSGw12+4hc
L8UN8o87+X00oXOeC74W8iPRp9P2xtahAQqrYov3aBgtG3K9LOvxGLvh4Gs/Q1T3
COagHohPM6+vOlzp414NSOd6glxiRLTCTgQdsBx14lwX4ZN0LZgxVXwpAsUBgN/X
OW8ZJCjK0Uh3y2tmOVNYQfQPHpWizpg4a/PioD6EX5B/AAySDiN6ktbb+nPBB0Q4
/BEamjE9v/V3/RLzOYQ9fKh/GY68Ocw7ine5dEsuErg2QQ1LWunM+aik5b08Jq0R
806wAX8zQandzgU21n23taNCfCWgCpWBLLMuUWJeUoUdHfUFEqz4B0qnJ9poaGFV
UzwZRHhMwkX3wD6yj2scf5jn1T1WLo/Ej6rPHMnEtODXXt8kJoqR8HHT/eCc83JE
8xTSBnjuZKnvXi1ZxeW01TXPVW+SrgAJv36jqvDxzCE7r+XBt4gZlUeX5I9qWJTp
YC6Eu0XQ+TNJHNcRVRcN6ozpbT+9du8013+/4Q8smWqjroM0H5O3p/VOYYxbUs+8
qIuVNF51sGFZA8Y1QwT++vB1pMNDthvWTFS/Qe3+bNjURruFOupgro85LkhmjVuG
qK40/GmLVkQq4Lhou7GcfsdsWmCduWBjdISJMxJp/irjNSDjxc5ucpBkFKzfZy1P
Zp9DahmvtNoAFpxNBlrJgUfq0Xp/JcyiSAAbcg5FRtEubkCoJwhemsfxROx0SAPA
/wmIk1Q6Rm4aXSXH/jTWr6K++dpPtNd9JI6Si57fJMVtG8MEhBMidmqGow+nHN/M
QWjhgxoaiY7DYGPeu3wDYLLwDhc13oTjmm3zNcnfbZuF8qG8RLld0T367csqlqRd
BYZP2Cxv3UjxJIOH4ImMumFwpwdq04zp8KnNf0s0dI2ntcQecWYyhX4p6vCMUvjo
ew5KEiKu1/AlO8I2NGLDCvVAXpoCHygPFPrUlZ5pRRoKd0pxA0gs/ldmlHHf4B1m
i+8pFHGpNi2vFs0VREvYBaD3JnejEMQVadcADUY6f1xMaR6SiIdnKjkmq89q9BfS
OEEsk6tGrxAejfD8aP8bAa+DIBycvfcqz0J+4LBzUhoUWadB22rs22yMX20o37qk
GMOCQ6So7QxADnGIMi7xPmyyyp645hvq/kuOXMiOp9B3bU27WkFNrda5j0bHnjKz
R7g1dhYQMhnSU4eK9SKS24TCjhHZgpX/m1IYkHOwFv6YXrU391QFog7y/AANi7Tz
jWFTdKXnQor/NTqLCjrFDusIqzI4zUdyle1WdU1zJTUgQe/kkb5HqTAQxO3E4Dem
jcKyEl/iNPyY2cIQq0YJRg==
//pragma protect end_data_block
//pragma protect digest_block
x7ApwIafMhdQyoSJ3LUp/7z63KI=
//pragma protect end_digest_block
//pragma protect end_protected
